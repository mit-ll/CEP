// File ./rom1.vhd translated with vhd2vl v2.4 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 1995

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002, 2005, 2008-2010 Larry Doolittle - LBNL
//     http://doolittle.icarus.com/~larry/vhd2vl/
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

// Rom file for twiddle factors 
// ../../../rtl/vhdl/WISHBONE_FFT/rom1.vhd contains 1024 points of 16 width 
//  for a 1024 point fft.
// no timescale needed

module rom1(
clk,
address,
datar,
datai
);

parameter [31:0] data_width=16;
parameter [31:0] address_width=10;
input clk;
input [9:0] address;
output [data_width - 1:0] datar;
output [data_width - 1:0] datai;

wire clk;
wire [9:0] address;
reg [data_width - 1:0] datar;
reg [data_width - 1:0] datai;
integer i;


  always @(posedge address or posedge clk) begin
    case(address)
    10'b 0000000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 0000000001 : begin
      datar <= 16'b 0111111111111101;
      datai <= 16'b 1111111001101110;
      //2
    end
    10'b 0000000010 : begin
      datar <= 16'b 0111111111110101;
      datai <= 16'b 1111110011011100;
      //4
    end
    10'b 0000000011 : begin
      datar <= 16'b 0111111111101001;
      datai <= 16'b 1111101101001010;
      //6
    end
    10'b 0000000100 : begin
      datar <= 16'b 0111111111011000;
      datai <= 16'b 1111100110111000;
      //8
    end
    10'b 0000000101 : begin
      datar <= 16'b 0111111111000001;
      datai <= 16'b 1111100000100111;
      //10
    end
    10'b 0000000110 : begin
      datar <= 16'b 0111111110100110;
      datai <= 16'b 1111011010010110;
      //12
    end
    10'b 0000000111 : begin
      datar <= 16'b 0111111110000110;
      datai <= 16'b 1111010100000101;
      //14
    end
    10'b 0000001000 : begin
      datar <= 16'b 0111111101100001;
      datai <= 16'b 1111001101110100;
      //16
    end
    10'b 0000001001 : begin
      datar <= 16'b 0111111100110111;
      datai <= 16'b 1111000111100100;
      //18
    end
    10'b 0000001010 : begin
      datar <= 16'b 0111111100001001;
      datai <= 16'b 1111000001010101;
      //20
    end
    10'b 0000001011 : begin
      datar <= 16'b 0111111011010101;
      datai <= 16'b 1110111011000110;
      //22
    end
    10'b 0000001100 : begin
      datar <= 16'b 0111111010011100;
      datai <= 16'b 1110110100111000;
      //24
    end
    10'b 0000001101 : begin
      datar <= 16'b 0111111001011111;
      datai <= 16'b 1110101110101011;
      //26
    end
    10'b 0000001110 : begin
      datar <= 16'b 0111111000011101;
      datai <= 16'b 1110101000011110;
      //28
    end
    10'b 0000001111 : begin
      datar <= 16'b 0111110111010101;
      datai <= 16'b 1110100010010010;
      //30
    end
    10'b 0000010000 : begin
      datar <= 16'b 0111110110001001;
      datai <= 16'b 1110011100000111;
      //32
    end
    10'b 0000010001 : begin
      datar <= 16'b 0111110100111001;
      datai <= 16'b 1110010101111110;
      //34
    end
    10'b 0000010010 : begin
      datar <= 16'b 0111110011100011;
      datai <= 16'b 1110001111110101;
      //36
    end
    10'b 0000010011 : begin
      datar <= 16'b 0111110010001000;
      datai <= 16'b 1110001001101101;
      //38
    end
    10'b 0000010100 : begin
      datar <= 16'b 0111110000101001;
      datai <= 16'b 1110000011100110;
      //40
    end
    10'b 0000010101 : begin
      datar <= 16'b 0111101111000101;
      datai <= 16'b 1101111101100001;
      //42
    end
    10'b 0000010110 : begin
      datar <= 16'b 0111101101011100;
      datai <= 16'b 1101110111011101;
      //44
    end
    10'b 0000010111 : begin
      datar <= 16'b 0111101011101110;
      datai <= 16'b 1101110001011010;
      //46
    end
    10'b 0000011000 : begin
      datar <= 16'b 0111101001111100;
      datai <= 16'b 1101101011011000;
      //48
    end
    10'b 0000011001 : begin
      datar <= 16'b 0111101000000101;
      datai <= 16'b 1101100101011000;
      //50
    end
    10'b 0000011010 : begin
      datar <= 16'b 0111100110001001;
      datai <= 16'b 1101011111011010;
      //52
    end
    10'b 0000011011 : begin
      datar <= 16'b 0111100100001001;
      datai <= 16'b 1101011001011101;
      //54
    end
    10'b 0000011100 : begin
      datar <= 16'b 0111100010000100;
      datai <= 16'b 1101010011100001;
      //56
    end
    10'b 0000011101 : begin
      datar <= 16'b 0111011111111010;
      datai <= 16'b 1101001101100111;
      //58
    end
    10'b 0000011110 : begin
      datar <= 16'b 0111011101101011;
      datai <= 16'b 1101000111101111;
      //60
    end
    10'b 0000011111 : begin
      datar <= 16'b 0111011011011000;
      datai <= 16'b 1101000001111001;
      //62
    end
    10'b 0000100000 : begin
      datar <= 16'b 0111011001000001;
      datai <= 16'b 1100111100000101;
      //64
    end
    10'b 0000100001 : begin
      datar <= 16'b 0111010110100101;
      datai <= 16'b 1100110110010010;
      //66
    end
    10'b 0000100010 : begin
      datar <= 16'b 0111010100000100;
      datai <= 16'b 1100110000100001;
      //68
    end
    10'b 0000100011 : begin
      datar <= 16'b 0111010001011111;
      datai <= 16'b 1100101010110011;
      //70
    end
    10'b 0000100100 : begin
      datar <= 16'b 0111001110110101;
      datai <= 16'b 1100100101000110;
      //72
    end
    10'b 0000100101 : begin
      datar <= 16'b 0111001100000111;
      datai <= 16'b 1100011111011100;
      //74
    end
    10'b 0000100110 : begin
      datar <= 16'b 0111001001010100;
      datai <= 16'b 1100011001110100;
      //76
    end
    10'b 0000100111 : begin
      datar <= 16'b 0111000110011101;
      datai <= 16'b 1100010100001110;
      //78
    end
    10'b 0000101000 : begin
      datar <= 16'b 0111000011100010;
      datai <= 16'b 1100001110101010;
      //80
    end
    10'b 0000101001 : begin
      datar <= 16'b 0111000000100010;
      datai <= 16'b 1100001001001000;
      //82
    end
    10'b 0000101010 : begin
      datar <= 16'b 0110111101011110;
      datai <= 16'b 1100000011101001;
      //84
    end
    10'b 0000101011 : begin
      datar <= 16'b 0110111010010110;
      datai <= 16'b 1011111110001101;
      //86
    end
    10'b 0000101100 : begin
      datar <= 16'b 0110110111001001;
      datai <= 16'b 1011111000110010;
      //88
    end
    10'b 0000101101 : begin
      datar <= 16'b 0110110011111000;
      datai <= 16'b 1011110011011011;
      //90
    end
    10'b 0000101110 : begin
      datar <= 16'b 0110110000100011;
      datai <= 16'b 1011101110000110;
      //92
    end
    10'b 0000101111 : begin
      datar <= 16'b 0110101101001010;
      datai <= 16'b 1011101000110011;
      //94
    end
    10'b 0000110000 : begin
      datar <= 16'b 0110101001101101;
      datai <= 16'b 1011100011100100;
      //96
    end
    10'b 0000110001 : begin
      datar <= 16'b 0110100110001011;
      datai <= 16'b 1011011110010111;
      //98
    end
    10'b 0000110010 : begin
      datar <= 16'b 0110100010100110;
      datai <= 16'b 1011011001001100;
      //100
    end
    10'b 0000110011 : begin
      datar <= 16'b 0110011110111100;
      datai <= 16'b 1011010100000101;
      //102
    end
    10'b 0000110100 : begin
      datar <= 16'b 0110011011001111;
      datai <= 16'b 1011001111000001;
      //104
    end
    10'b 0000110101 : begin
      datar <= 16'b 0110010111011101;
      datai <= 16'b 1011001001111111;
      //106
    end
    10'b 0000110110 : begin
      datar <= 16'b 0110010011101000;
      datai <= 16'b 1011000101000001;
      //108
    end
    10'b 0000110111 : begin
      datar <= 16'b 0110001111101110;
      datai <= 16'b 1011000000000101;
      //110
    end
    10'b 0000111000 : begin
      datar <= 16'b 0110001011110001;
      datai <= 16'b 1010111011001101;
      //112
    end
    10'b 0000111001 : begin
      datar <= 16'b 0110000111110000;
      datai <= 16'b 1010110110011000;
      //114
    end
    10'b 0000111010 : begin
      datar <= 16'b 0110000011101011;
      datai <= 16'b 1010110001100101;
      //116
    end
    10'b 0000111011 : begin
      datar <= 16'b 0101111111100011;
      datai <= 16'b 1010101100110111;
      //118
    end
    10'b 0000111100 : begin
      datar <= 16'b 0101111011010111;
      datai <= 16'b 1010101000001011;
      //120
    end
    10'b 0000111101 : begin
      datar <= 16'b 0101110111000111;
      datai <= 16'b 1010100011100011;
      //122
    end
    10'b 0000111110 : begin
      datar <= 16'b 0101110010110011;
      datai <= 16'b 1010011110111110;
      //124
    end
    10'b 0000111111 : begin
      datar <= 16'b 0101101110011100;
      datai <= 16'b 1010011010011100;
      //126
    end
    10'b 0001000000 : begin
      datar <= 16'b 0101101010000010;
      datai <= 16'b 1010010101111110;
      //128
    end
    10'b 0001000001 : begin
      datar <= 16'b 0101100101100100;
      datai <= 16'b 1010010001100100;
      //130
    end
    10'b 0001000010 : begin
      datar <= 16'b 0101100001000010;
      datai <= 16'b 1010001101001101;
      //132
    end
    10'b 0001000011 : begin
      datar <= 16'b 0101011100011101;
      datai <= 16'b 1010001000111001;
      //134
    end
    10'b 0001000100 : begin
      datar <= 16'b 0101010111110101;
      datai <= 16'b 1010000100101001;
      //136
    end
    10'b 0001000101 : begin
      datar <= 16'b 0101010011001001;
      datai <= 16'b 1010000000011101;
      //138
    end
    10'b 0001000110 : begin
      datar <= 16'b 0101001110011011;
      datai <= 16'b 1001111100010101;
      //140
    end
    10'b 0001000111 : begin
      datar <= 16'b 0101001001101000;
      datai <= 16'b 1001111000010000;
      //142
    end
    10'b 0001001000 : begin
      datar <= 16'b 0101000100110011;
      datai <= 16'b 1001110100001111;
      //144
    end
    10'b 0001001001 : begin
      datar <= 16'b 0100111111111011;
      datai <= 16'b 1001110000010010;
      //146
    end
    10'b 0001001010 : begin
      datar <= 16'b 0100111010111111;
      datai <= 16'b 1001101100011000;
      //148
    end
    10'b 0001001011 : begin
      datar <= 16'b 0100110110000001;
      datai <= 16'b 1001101000100011;
      //150
    end
    10'b 0001001100 : begin
      datar <= 16'b 0100110000111111;
      datai <= 16'b 1001100100110001;
      //152
    end
    10'b 0001001101 : begin
      datar <= 16'b 0100101011111011;
      datai <= 16'b 1001100001000100;
      //154
    end
    10'b 0001001110 : begin
      datar <= 16'b 0100100110110100;
      datai <= 16'b 1001011101011010;
      //156
    end
    10'b 0001001111 : begin
      datar <= 16'b 0100100001101001;
      datai <= 16'b 1001011001110101;
      //158
    end
    10'b 0001010000 : begin
      datar <= 16'b 0100011100011100;
      datai <= 16'b 1001010110010011;
      //160
    end
    10'b 0001010001 : begin
      datar <= 16'b 0100010111001101;
      datai <= 16'b 1001010010110110;
      //162
    end
    10'b 0001010010 : begin
      datar <= 16'b 0100010001111010;
      datai <= 16'b 1001001111011101;
      //164
    end
    10'b 0001010011 : begin
      datar <= 16'b 0100001100100101;
      datai <= 16'b 1001001100001000;
      //166
    end
    10'b 0001010100 : begin
      datar <= 16'b 0100000111001110;
      datai <= 16'b 1001001000110111;
      //168
    end
    10'b 0001010101 : begin
      datar <= 16'b 0100000001110011;
      datai <= 16'b 1001000101101010;
      //170
    end
    10'b 0001010110 : begin
      datar <= 16'b 0011111100010111;
      datai <= 16'b 1001000010100010;
      //172
    end
    10'b 0001010111 : begin
      datar <= 16'b 0011110110111000;
      datai <= 16'b 1000111111011110;
      //174
    end
    10'b 0001011000 : begin
      datar <= 16'b 0011110001010110;
      datai <= 16'b 1000111100011110;
      //176
    end
    10'b 0001011001 : begin
      datar <= 16'b 0011101011110010;
      datai <= 16'b 1000111001100011;
      //178
    end
    10'b 0001011010 : begin
      datar <= 16'b 0011100110001100;
      datai <= 16'b 1000110110101100;
      //180
    end
    10'b 0001011011 : begin
      datar <= 16'b 0011100000100100;
      datai <= 16'b 1000110011111001;
      //182
    end
    10'b 0001011100 : begin
      datar <= 16'b 0011011010111010;
      datai <= 16'b 1000110001001011;
      //184
    end
    10'b 0001011101 : begin
      datar <= 16'b 0011010101001101;
      datai <= 16'b 1000101110100001;
      //186
    end
    10'b 0001011110 : begin
      datar <= 16'b 0011001111011111;
      datai <= 16'b 1000101011111100;
      //188
    end
    10'b 0001011111 : begin
      datar <= 16'b 0011001001101110;
      datai <= 16'b 1000101001011011;
      //190
    end
    10'b 0001100000 : begin
      datar <= 16'b 0011000011111011;
      datai <= 16'b 1000100110111111;
      //192
    end
    10'b 0001100001 : begin
      datar <= 16'b 0010111110000111;
      datai <= 16'b 1000100100101000;
      //194
    end
    10'b 0001100010 : begin
      datar <= 16'b 0010111000010001;
      datai <= 16'b 1000100010010101;
      //196
    end
    10'b 0001100011 : begin
      datar <= 16'b 0010110010011001;
      datai <= 16'b 1000100000000110;
      //198
    end
    10'b 0001100100 : begin
      datar <= 16'b 0010101100011111;
      datai <= 16'b 1000011101111100;
      //200
    end
    10'b 0001100101 : begin
      datar <= 16'b 0010100110100011;
      datai <= 16'b 1000011011110111;
      //202
    end
    10'b 0001100110 : begin
      datar <= 16'b 0010100000100110;
      datai <= 16'b 1000011001110111;
      //204
    end
    10'b 0001100111 : begin
      datar <= 16'b 0010011010101000;
      datai <= 16'b 1000010111111011;
      //206
    end
    10'b 0001101000 : begin
      datar <= 16'b 0010010100101000;
      datai <= 16'b 1000010110000100;
      //208
    end
    10'b 0001101001 : begin
      datar <= 16'b 0010001110100110;
      datai <= 16'b 1000010100010010;
      //210
    end
    10'b 0001101010 : begin
      datar <= 16'b 0010001000100011;
      datai <= 16'b 1000010010100100;
      //212
    end
    10'b 0001101011 : begin
      datar <= 16'b 0010000010011111;
      datai <= 16'b 1000010000111011;
      //214
    end
    10'b 0001101100 : begin
      datar <= 16'b 0001111100011010;
      datai <= 16'b 1000001111010111;
      //216
    end
    10'b 0001101101 : begin
      datar <= 16'b 0001110110010011;
      datai <= 16'b 1000001101111000;
      //218
    end
    10'b 0001101110 : begin
      datar <= 16'b 0001110000001011;
      datai <= 16'b 1000001100011101;
      //220
    end
    10'b 0001101111 : begin
      datar <= 16'b 0001101010000010;
      datai <= 16'b 1000001011000111;
      //222
    end
    10'b 0001110000 : begin
      datar <= 16'b 0001100011111001;
      datai <= 16'b 1000001001110111;
      //224
    end
    10'b 0001110001 : begin
      datar <= 16'b 0001011101101110;
      datai <= 16'b 1000001000101011;
      //226
    end
    10'b 0001110010 : begin
      datar <= 16'b 0001010111100010;
      datai <= 16'b 1000000111100011;
      //228
    end
    10'b 0001110011 : begin
      datar <= 16'b 0001010001010101;
      datai <= 16'b 1000000110100001;
      //230
    end
    10'b 0001110100 : begin
      datar <= 16'b 0001001011001000;
      datai <= 16'b 1000000101100100;
      //232
    end
    10'b 0001110101 : begin
      datar <= 16'b 0001000100111010;
      datai <= 16'b 1000000100101011;
      //234
    end
    10'b 0001110110 : begin
      datar <= 16'b 0000111110101011;
      datai <= 16'b 1000000011110111;
      //236
    end
    10'b 0001110111 : begin
      datar <= 16'b 0000111000011100;
      datai <= 16'b 1000000011001001;
      //238
    end
    10'b 0001111000 : begin
      datar <= 16'b 0000110010001100;
      datai <= 16'b 1000000010011111;
      //240
    end
    10'b 0001111001 : begin
      datar <= 16'b 0000101011111011;
      datai <= 16'b 1000000001111010;
      //242
    end
    10'b 0001111010 : begin
      datar <= 16'b 0000100101101010;
      datai <= 16'b 1000000001011010;
      //244
    end
    10'b 0001111011 : begin
      datar <= 16'b 0000011111011001;
      datai <= 16'b 1000000000111111;
      //246
    end
    10'b 0001111100 : begin
      datar <= 16'b 0000011001001000;
      datai <= 16'b 1000000000101000;
      //248
    end
    10'b 0001111101 : begin
      datar <= 16'b 0000010010110110;
      datai <= 16'b 1000000000010111;
      //250
    end
    10'b 0001111110 : begin
      datar <= 16'b 0000001100100100;
      datai <= 16'b 1000000000001011;
      //252
    end
    10'b 0001111111 : begin
      datar <= 16'b 0000000110010010;
      datai <= 16'b 1000000000000011;
      //254
    end
    10'b 0010000000 : begin
      datar <= 16'b 0000000000000000;
      datai <= 16'b 1000000000000001;
      //256
    end
    10'b 0010000001 : begin
      datar <= 16'b 1111111001101110;
      datai <= 16'b 1000000000000011;
      //258
    end
    10'b 0010000010 : begin
      datar <= 16'b 1111110011011100;
      datai <= 16'b 1000000000001011;
      //260
    end
    10'b 0010000011 : begin
      datar <= 16'b 1111101101001010;
      datai <= 16'b 1000000000010111;
      //262
    end
    10'b 0010000100 : begin
      datar <= 16'b 1111100110111000;
      datai <= 16'b 1000000000101000;
      //264
    end
    10'b 0010000101 : begin
      datar <= 16'b 1111100000100111;
      datai <= 16'b 1000000000111111;
      //266
    end
    10'b 0010000110 : begin
      datar <= 16'b 1111011010010110;
      datai <= 16'b 1000000001011010;
      //268
    end
    10'b 0010000111 : begin
      datar <= 16'b 1111010100000101;
      datai <= 16'b 1000000001111010;
      //270
    end
    10'b 0010001000 : begin
      datar <= 16'b 1111001101110100;
      datai <= 16'b 1000000010011111;
      //272
    end
    10'b 0010001001 : begin
      datar <= 16'b 1111000111100100;
      datai <= 16'b 1000000011001001;
      //274
    end
    10'b 0010001010 : begin
      datar <= 16'b 1111000001010101;
      datai <= 16'b 1000000011110111;
      //276
    end
    10'b 0010001011 : begin
      datar <= 16'b 1110111011000110;
      datai <= 16'b 1000000100101011;
      //278
    end
    10'b 0010001100 : begin
      datar <= 16'b 1110110100111000;
      datai <= 16'b 1000000101100100;
      //280
    end
    10'b 0010001101 : begin
      datar <= 16'b 1110101110101011;
      datai <= 16'b 1000000110100001;
      //282
    end
    10'b 0010001110 : begin
      datar <= 16'b 1110101000011110;
      datai <= 16'b 1000000111100011;
      //284
    end
    10'b 0010001111 : begin
      datar <= 16'b 1110100010010010;
      datai <= 16'b 1000001000101011;
      //286
    end
    10'b 0010010000 : begin
      datar <= 16'b 1110011100000111;
      datai <= 16'b 1000001001110111;
      //288
    end
    10'b 0010010001 : begin
      datar <= 16'b 1110010101111110;
      datai <= 16'b 1000001011000111;
      //290
    end
    10'b 0010010010 : begin
      datar <= 16'b 1110001111110101;
      datai <= 16'b 1000001100011101;
      //292
    end
    10'b 0010010011 : begin
      datar <= 16'b 1110001001101101;
      datai <= 16'b 1000001101111000;
      //294
    end
    10'b 0010010100 : begin
      datar <= 16'b 1110000011100110;
      datai <= 16'b 1000001111010111;
      //296
    end
    10'b 0010010101 : begin
      datar <= 16'b 1101111101100001;
      datai <= 16'b 1000010000111011;
      //298
    end
    10'b 0010010110 : begin
      datar <= 16'b 1101110111011101;
      datai <= 16'b 1000010010100100;
      //300
    end
    10'b 0010010111 : begin
      datar <= 16'b 1101110001011010;
      datai <= 16'b 1000010100010010;
      //302
    end
    10'b 0010011000 : begin
      datar <= 16'b 1101101011011000;
      datai <= 16'b 1000010110000100;
      //304
    end
    10'b 0010011001 : begin
      datar <= 16'b 1101100101011000;
      datai <= 16'b 1000010111111011;
      //306
    end
    10'b 0010011010 : begin
      datar <= 16'b 1101011111011010;
      datai <= 16'b 1000011001110111;
      //308
    end
    10'b 0010011011 : begin
      datar <= 16'b 1101011001011101;
      datai <= 16'b 1000011011110111;
      //310
    end
    10'b 0010011100 : begin
      datar <= 16'b 1101010011100001;
      datai <= 16'b 1000011101111100;
      //312
    end
    10'b 0010011101 : begin
      datar <= 16'b 1101001101100111;
      datai <= 16'b 1000100000000110;
      //314
    end
    10'b 0010011110 : begin
      datar <= 16'b 1101000111101111;
      datai <= 16'b 1000100010010101;
      //316
    end
    10'b 0010011111 : begin
      datar <= 16'b 1101000001111001;
      datai <= 16'b 1000100100101000;
      //318
    end
    10'b 0010100000 : begin
      datar <= 16'b 1100111100000101;
      datai <= 16'b 1000100110111111;
      //320
    end
    10'b 0010100001 : begin
      datar <= 16'b 1100110110010010;
      datai <= 16'b 1000101001011011;
      //322
    end
    10'b 0010100010 : begin
      datar <= 16'b 1100110000100001;
      datai <= 16'b 1000101011111100;
      //324
    end
    10'b 0010100011 : begin
      datar <= 16'b 1100101010110011;
      datai <= 16'b 1000101110100001;
      //326
    end
    10'b 0010100100 : begin
      datar <= 16'b 1100100101000110;
      datai <= 16'b 1000110001001011;
      //328
    end
    10'b 0010100101 : begin
      datar <= 16'b 1100011111011100;
      datai <= 16'b 1000110011111001;
      //330
    end
    10'b 0010100110 : begin
      datar <= 16'b 1100011001110100;
      datai <= 16'b 1000110110101100;
      //332
    end
    10'b 0010100111 : begin
      datar <= 16'b 1100010100001110;
      datai <= 16'b 1000111001100011;
      //334
    end
    10'b 0010101000 : begin
      datar <= 16'b 1100001110101010;
      datai <= 16'b 1000111100011110;
      //336
    end
    10'b 0010101001 : begin
      datar <= 16'b 1100001001001000;
      datai <= 16'b 1000111111011110;
      //338
    end
    10'b 0010101010 : begin
      datar <= 16'b 1100000011101001;
      datai <= 16'b 1001000010100010;
      //340
    end
    10'b 0010101011 : begin
      datar <= 16'b 1011111110001101;
      datai <= 16'b 1001000101101010;
      //342
    end
    10'b 0010101100 : begin
      datar <= 16'b 1011111000110010;
      datai <= 16'b 1001001000110111;
      //344
    end
    10'b 0010101101 : begin
      datar <= 16'b 1011110011011011;
      datai <= 16'b 1001001100001000;
      //346
    end
    10'b 0010101110 : begin
      datar <= 16'b 1011101110000110;
      datai <= 16'b 1001001111011101;
      //348
    end
    10'b 0010101111 : begin
      datar <= 16'b 1011101000110011;
      datai <= 16'b 1001010010110110;
      //350
    end
    10'b 0010110000 : begin
      datar <= 16'b 1011100011100100;
      datai <= 16'b 1001010110010011;
      //352
    end
    10'b 0010110001 : begin
      datar <= 16'b 1011011110010111;
      datai <= 16'b 1001011001110101;
      //354
    end
    10'b 0010110010 : begin
      datar <= 16'b 1011011001001100;
      datai <= 16'b 1001011101011010;
      //356
    end
    10'b 0010110011 : begin
      datar <= 16'b 1011010100000101;
      datai <= 16'b 1001100001000100;
      //358
    end
    10'b 0010110100 : begin
      datar <= 16'b 1011001111000001;
      datai <= 16'b 1001100100110001;
      //360
    end
    10'b 0010110101 : begin
      datar <= 16'b 1011001001111111;
      datai <= 16'b 1001101000100011;
      //362
    end
    10'b 0010110110 : begin
      datar <= 16'b 1011000101000001;
      datai <= 16'b 1001101100011000;
      //364
    end
    10'b 0010110111 : begin
      datar <= 16'b 1011000000000101;
      datai <= 16'b 1001110000010010;
      //366
    end
    10'b 0010111000 : begin
      datar <= 16'b 1010111011001101;
      datai <= 16'b 1001110100001111;
      //368
    end
    10'b 0010111001 : begin
      datar <= 16'b 1010110110011000;
      datai <= 16'b 1001111000010000;
      //370
    end
    10'b 0010111010 : begin
      datar <= 16'b 1010110001100101;
      datai <= 16'b 1001111100010101;
      //372
    end
    10'b 0010111011 : begin
      datar <= 16'b 1010101100110111;
      datai <= 16'b 1010000000011101;
      //374
    end
    10'b 0010111100 : begin
      datar <= 16'b 1010101000001011;
      datai <= 16'b 1010000100101001;
      //376
    end
    10'b 0010111101 : begin
      datar <= 16'b 1010100011100011;
      datai <= 16'b 1010001000111001;
      //378
    end
    10'b 0010111110 : begin
      datar <= 16'b 1010011110111110;
      datai <= 16'b 1010001101001101;
      //380
    end
    10'b 0010111111 : begin
      datar <= 16'b 1010011010011100;
      datai <= 16'b 1010010001100100;
      //382
    end
    10'b 0011000000 : begin
      datar <= 16'b 1010010101111110;
      datai <= 16'b 1010010101111110;
      //384
    end
    10'b 0011000001 : begin
      datar <= 16'b 1010010001100100;
      datai <= 16'b 1010011010011100;
      //386
    end
    10'b 0011000010 : begin
      datar <= 16'b 1010001101001101;
      datai <= 16'b 1010011110111110;
      //388
    end
    10'b 0011000011 : begin
      datar <= 16'b 1010001000111001;
      datai <= 16'b 1010100011100011;
      //390
    end
    10'b 0011000100 : begin
      datar <= 16'b 1010000100101001;
      datai <= 16'b 1010101000001011;
      //392
    end
    10'b 0011000101 : begin
      datar <= 16'b 1010000000011101;
      datai <= 16'b 1010101100110111;
      //394
    end
    10'b 0011000110 : begin
      datar <= 16'b 1001111100010101;
      datai <= 16'b 1010110001100101;
      //396
    end
    10'b 0011000111 : begin
      datar <= 16'b 1001111000010000;
      datai <= 16'b 1010110110011000;
      //398
    end
    10'b 0011001000 : begin
      datar <= 16'b 1001110100001111;
      datai <= 16'b 1010111011001101;
      //400
    end
    10'b 0011001001 : begin
      datar <= 16'b 1001110000010010;
      datai <= 16'b 1011000000000101;
      //402
    end
    10'b 0011001010 : begin
      datar <= 16'b 1001101100011000;
      datai <= 16'b 1011000101000001;
      //404
    end
    10'b 0011001011 : begin
      datar <= 16'b 1001101000100011;
      datai <= 16'b 1011001001111111;
      //406
    end
    10'b 0011001100 : begin
      datar <= 16'b 1001100100110001;
      datai <= 16'b 1011001111000001;
      //408
    end
    10'b 0011001101 : begin
      datar <= 16'b 1001100001000100;
      datai <= 16'b 1011010100000101;
      //410
    end
    10'b 0011001110 : begin
      datar <= 16'b 1001011101011010;
      datai <= 16'b 1011011001001100;
      //412
    end
    10'b 0011001111 : begin
      datar <= 16'b 1001011001110101;
      datai <= 16'b 1011011110010111;
      //414
    end
    10'b 0011010000 : begin
      datar <= 16'b 1001010110010011;
      datai <= 16'b 1011100011100100;
      //416
    end
    10'b 0011010001 : begin
      datar <= 16'b 1001010010110110;
      datai <= 16'b 1011101000110011;
      //418
    end
    10'b 0011010010 : begin
      datar <= 16'b 1001001111011101;
      datai <= 16'b 1011101110000110;
      //420
    end
    10'b 0011010011 : begin
      datar <= 16'b 1001001100001000;
      datai <= 16'b 1011110011011011;
      //422
    end
    10'b 0011010100 : begin
      datar <= 16'b 1001001000110111;
      datai <= 16'b 1011111000110010;
      //424
    end
    10'b 0011010101 : begin
      datar <= 16'b 1001000101101010;
      datai <= 16'b 1011111110001101;
      //426
    end
    10'b 0011010110 : begin
      datar <= 16'b 1001000010100010;
      datai <= 16'b 1100000011101001;
      //428
    end
    10'b 0011010111 : begin
      datar <= 16'b 1000111111011110;
      datai <= 16'b 1100001001001000;
      //430
    end
    10'b 0011011000 : begin
      datar <= 16'b 1000111100011110;
      datai <= 16'b 1100001110101010;
      //432
    end
    10'b 0011011001 : begin
      datar <= 16'b 1000111001100011;
      datai <= 16'b 1100010100001110;
      //434
    end
    10'b 0011011010 : begin
      datar <= 16'b 1000110110101100;
      datai <= 16'b 1100011001110100;
      //436
    end
    10'b 0011011011 : begin
      datar <= 16'b 1000110011111001;
      datai <= 16'b 1100011111011100;
      //438
    end
    10'b 0011011100 : begin
      datar <= 16'b 1000110001001011;
      datai <= 16'b 1100100101000110;
      //440
    end
    10'b 0011011101 : begin
      datar <= 16'b 1000101110100001;
      datai <= 16'b 1100101010110011;
      //442
    end
    10'b 0011011110 : begin
      datar <= 16'b 1000101011111100;
      datai <= 16'b 1100110000100001;
      //444
    end
    10'b 0011011111 : begin
      datar <= 16'b 1000101001011011;
      datai <= 16'b 1100110110010010;
      //446
    end
    10'b 0011100000 : begin
      datar <= 16'b 1000100110111111;
      datai <= 16'b 1100111100000101;
      //448
    end
    10'b 0011100001 : begin
      datar <= 16'b 1000100100101000;
      datai <= 16'b 1101000001111001;
      //450
    end
    10'b 0011100010 : begin
      datar <= 16'b 1000100010010101;
      datai <= 16'b 1101000111101111;
      //452
    end
    10'b 0011100011 : begin
      datar <= 16'b 1000100000000110;
      datai <= 16'b 1101001101100111;
      //454
    end
    10'b 0011100100 : begin
      datar <= 16'b 1000011101111100;
      datai <= 16'b 1101010011100001;
      //456
    end
    10'b 0011100101 : begin
      datar <= 16'b 1000011011110111;
      datai <= 16'b 1101011001011101;
      //458
    end
    10'b 0011100110 : begin
      datar <= 16'b 1000011001110111;
      datai <= 16'b 1101011111011010;
      //460
    end
    10'b 0011100111 : begin
      datar <= 16'b 1000010111111011;
      datai <= 16'b 1101100101011000;
      //462
    end
    10'b 0011101000 : begin
      datar <= 16'b 1000010110000100;
      datai <= 16'b 1101101011011000;
      //464
    end
    10'b 0011101001 : begin
      datar <= 16'b 1000010100010010;
      datai <= 16'b 1101110001011010;
      //466
    end
    10'b 0011101010 : begin
      datar <= 16'b 1000010010100100;
      datai <= 16'b 1101110111011101;
      //468
    end
    10'b 0011101011 : begin
      datar <= 16'b 1000010000111011;
      datai <= 16'b 1101111101100001;
      //470
    end
    10'b 0011101100 : begin
      datar <= 16'b 1000001111010111;
      datai <= 16'b 1110000011100110;
      //472
    end
    10'b 0011101101 : begin
      datar <= 16'b 1000001101111000;
      datai <= 16'b 1110001001101101;
      //474
    end
    10'b 0011101110 : begin
      datar <= 16'b 1000001100011101;
      datai <= 16'b 1110001111110101;
      //476
    end
    10'b 0011101111 : begin
      datar <= 16'b 1000001011000111;
      datai <= 16'b 1110010101111110;
      //478
    end
    10'b 0011110000 : begin
      datar <= 16'b 1000001001110111;
      datai <= 16'b 1110011100000111;
      //480
    end
    10'b 0011110001 : begin
      datar <= 16'b 1000001000101011;
      datai <= 16'b 1110100010010010;
      //482
    end
    10'b 0011110010 : begin
      datar <= 16'b 1000000111100011;
      datai <= 16'b 1110101000011110;
      //484
    end
    10'b 0011110011 : begin
      datar <= 16'b 1000000110100001;
      datai <= 16'b 1110101110101011;
      //486
    end
    10'b 0011110100 : begin
      datar <= 16'b 1000000101100100;
      datai <= 16'b 1110110100111000;
      //488
    end
    10'b 0011110101 : begin
      datar <= 16'b 1000000100101011;
      datai <= 16'b 1110111011000110;
      //490
    end
    10'b 0011110110 : begin
      datar <= 16'b 1000000011110111;
      datai <= 16'b 1111000001010101;
      //492
    end
    10'b 0011110111 : begin
      datar <= 16'b 1000000011001001;
      datai <= 16'b 1111000111100100;
      //494
    end
    10'b 0011111000 : begin
      datar <= 16'b 1000000010011111;
      datai <= 16'b 1111001101110100;
      //496
    end
    10'b 0011111001 : begin
      datar <= 16'b 1000000001111010;
      datai <= 16'b 1111010100000101;
      //498
    end
    10'b 0011111010 : begin
      datar <= 16'b 1000000001011010;
      datai <= 16'b 1111011010010110;
      //500
    end
    10'b 0011111011 : begin
      datar <= 16'b 1000000000111111;
      datai <= 16'b 1111100000100111;
      //502
    end
    10'b 0011111100 : begin
      datar <= 16'b 1000000000101000;
      datai <= 16'b 1111100110111000;
      //504
    end
    10'b 0011111101 : begin
      datar <= 16'b 1000000000010111;
      datai <= 16'b 1111101101001010;
      //506
    end
    10'b 0011111110 : begin
      datar <= 16'b 1000000000001011;
      datai <= 16'b 1111110011011100;
      //508
    end
    10'b 0011111111 : begin
      datar <= 16'b 1000000000000011;
      datai <= 16'b 1111111001101110;
      //510
    end
    10'b 0100000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 0100000001 : begin
      datar <= 16'b 0111111111111110;
      datai <= 16'b 1111111100110111;
      //1
    end
    10'b 0100000010 : begin
      datar <= 16'b 0111111111111101;
      datai <= 16'b 1111111001101110;
      //2
    end
    10'b 0100000011 : begin
      datar <= 16'b 0111111111111001;
      datai <= 16'b 1111110110100101;
      //3
    end
    10'b 0100000100 : begin
      datar <= 16'b 0111111111110101;
      datai <= 16'b 1111110011011100;
      //4
    end
    10'b 0100000101 : begin
      datar <= 16'b 0111111111110000;
      datai <= 16'b 1111110000010011;
      //5
    end
    10'b 0100000110 : begin
      datar <= 16'b 0111111111101001;
      datai <= 16'b 1111101101001010;
      //6
    end
    10'b 0100000111 : begin
      datar <= 16'b 0111111111100001;
      datai <= 16'b 1111101010000001;
      //7
    end
    10'b 0100001000 : begin
      datar <= 16'b 0111111111011000;
      datai <= 16'b 1111100110111000;
      //8
    end
    10'b 0100001001 : begin
      datar <= 16'b 0111111111001101;
      datai <= 16'b 1111100011101111;
      //9
    end
    10'b 0100001010 : begin
      datar <= 16'b 0111111111000001;
      datai <= 16'b 1111100000100111;
      //10
    end
    10'b 0100001011 : begin
      datar <= 16'b 0111111110110100;
      datai <= 16'b 1111011101011110;
      //11
    end
    10'b 0100001100 : begin
      datar <= 16'b 0111111110100110;
      datai <= 16'b 1111011010010110;
      //12
    end
    10'b 0100001101 : begin
      datar <= 16'b 0111111110010111;
      datai <= 16'b 1111010111001101;
      //13
    end
    10'b 0100001110 : begin
      datar <= 16'b 0111111110000110;
      datai <= 16'b 1111010100000101;
      //14
    end
    10'b 0100001111 : begin
      datar <= 16'b 0111111101110100;
      datai <= 16'b 1111010000111100;
      //15
    end
    10'b 0100010000 : begin
      datar <= 16'b 0111111101100001;
      datai <= 16'b 1111001101110100;
      //16
    end
    10'b 0100010001 : begin
      datar <= 16'b 0111111101001101;
      datai <= 16'b 1111001010101100;
      //17
    end
    10'b 0100010010 : begin
      datar <= 16'b 0111111100110111;
      datai <= 16'b 1111000111100100;
      //18
    end
    10'b 0100010011 : begin
      datar <= 16'b 0111111100100001;
      datai <= 16'b 1111000100011101;
      //19
    end
    10'b 0100010100 : begin
      datar <= 16'b 0111111100001001;
      datai <= 16'b 1111000001010101;
      //20
    end
    10'b 0100010101 : begin
      datar <= 16'b 0111111011101111;
      datai <= 16'b 1110111110001110;
      //21
    end
    10'b 0100010110 : begin
      datar <= 16'b 0111111011010101;
      datai <= 16'b 1110111011000110;
      //22
    end
    10'b 0100010111 : begin
      datar <= 16'b 0111111010111001;
      datai <= 16'b 1110110111111111;
      //23
    end
    10'b 0100011000 : begin
      datar <= 16'b 0111111010011100;
      datai <= 16'b 1110110100111000;
      //24
    end
    10'b 0100011001 : begin
      datar <= 16'b 0111111001111110;
      datai <= 16'b 1110110001110001;
      //25
    end
    10'b 0100011010 : begin
      datar <= 16'b 0111111001011111;
      datai <= 16'b 1110101110101011;
      //26
    end
    10'b 0100011011 : begin
      datar <= 16'b 0111111000111110;
      datai <= 16'b 1110101011100100;
      //27
    end
    10'b 0100011100 : begin
      datar <= 16'b 0111111000011101;
      datai <= 16'b 1110101000011110;
      //28
    end
    10'b 0100011101 : begin
      datar <= 16'b 0111110111111010;
      datai <= 16'b 1110100101011000;
      //29
    end
    10'b 0100011110 : begin
      datar <= 16'b 0111110111010101;
      datai <= 16'b 1110100010010010;
      //30
    end
    10'b 0100011111 : begin
      datar <= 16'b 0111110110110000;
      datai <= 16'b 1110011111001101;
      //31
    end
    10'b 0100100000 : begin
      datar <= 16'b 0111110110001001;
      datai <= 16'b 1110011100000111;
      //32
    end
    10'b 0100100001 : begin
      datar <= 16'b 0111110101100010;
      datai <= 16'b 1110011001000010;
      //33
    end
    10'b 0100100010 : begin
      datar <= 16'b 0111110100111001;
      datai <= 16'b 1110010101111110;
      //34
    end
    10'b 0100100011 : begin
      datar <= 16'b 0111110100001110;
      datai <= 16'b 1110010010111001;
      //35
    end
    10'b 0100100100 : begin
      datar <= 16'b 0111110011100011;
      datai <= 16'b 1110001111110101;
      //36
    end
    10'b 0100100101 : begin
      datar <= 16'b 0111110010110110;
      datai <= 16'b 1110001100110001;
      //37
    end
    10'b 0100100110 : begin
      datar <= 16'b 0111110010001000;
      datai <= 16'b 1110001001101101;
      //38
    end
    10'b 0100100111 : begin
      datar <= 16'b 0111110001011001;
      datai <= 16'b 1110000110101001;
      //39
    end
    10'b 0100101000 : begin
      datar <= 16'b 0111110000101001;
      datai <= 16'b 1110000011100110;
      //40
    end
    10'b 0100101001 : begin
      datar <= 16'b 0111101111111000;
      datai <= 16'b 1110000000100011;
      //41
    end
    10'b 0100101010 : begin
      datar <= 16'b 0111101111000101;
      datai <= 16'b 1101111101100001;
      //42
    end
    10'b 0100101011 : begin
      datar <= 16'b 0111101110010001;
      datai <= 16'b 1101111010011111;
      //43
    end
    10'b 0100101100 : begin
      datar <= 16'b 0111101101011100;
      datai <= 16'b 1101110111011101;
      //44
    end
    10'b 0100101101 : begin
      datar <= 16'b 0111101100100110;
      datai <= 16'b 1101110100011011;
      //45
    end
    10'b 0100101110 : begin
      datar <= 16'b 0111101011101110;
      datai <= 16'b 1101110001011010;
      //46
    end
    10'b 0100101111 : begin
      datar <= 16'b 0111101010110110;
      datai <= 16'b 1101101110011001;
      //47
    end
    10'b 0100110000 : begin
      datar <= 16'b 0111101001111100;
      datai <= 16'b 1101101011011000;
      //48
    end
    10'b 0100110001 : begin
      datar <= 16'b 0111101001000001;
      datai <= 16'b 1101101000011000;
      //49
    end
    10'b 0100110010 : begin
      datar <= 16'b 0111101000000101;
      datai <= 16'b 1101100101011000;
      //50
    end
    10'b 0100110011 : begin
      datar <= 16'b 0111100111001000;
      datai <= 16'b 1101100010011001;
      //51
    end
    10'b 0100110100 : begin
      datar <= 16'b 0111100110001001;
      datai <= 16'b 1101011111011010;
      //52
    end
    10'b 0100110101 : begin
      datar <= 16'b 0111100101001010;
      datai <= 16'b 1101011100011011;
      //53
    end
    10'b 0100110110 : begin
      datar <= 16'b 0111100100001001;
      datai <= 16'b 1101011001011101;
      //54
    end
    10'b 0100110111 : begin
      datar <= 16'b 0111100011000111;
      datai <= 16'b 1101010110011111;
      //55
    end
    10'b 0100111000 : begin
      datar <= 16'b 0111100010000100;
      datai <= 16'b 1101010011100001;
      //56
    end
    10'b 0100111001 : begin
      datar <= 16'b 0111100000111111;
      datai <= 16'b 1101010000100100;
      //57
    end
    10'b 0100111010 : begin
      datar <= 16'b 0111011111111010;
      datai <= 16'b 1101001101100111;
      //58
    end
    10'b 0100111011 : begin
      datar <= 16'b 0111011110110011;
      datai <= 16'b 1101001010101011;
      //59
    end
    10'b 0100111100 : begin
      datar <= 16'b 0111011101101011;
      datai <= 16'b 1101000111101111;
      //60
    end
    10'b 0100111101 : begin
      datar <= 16'b 0111011100100010;
      datai <= 16'b 1101000100110100;
      //61
    end
    10'b 0100111110 : begin
      datar <= 16'b 0111011011011000;
      datai <= 16'b 1101000001111001;
      //62
    end
    10'b 0100111111 : begin
      datar <= 16'b 0111011010001101;
      datai <= 16'b 1100111110111111;
      //63
    end
    10'b 0101000000 : begin
      datar <= 16'b 0111011001000001;
      datai <= 16'b 1100111100000101;
      //64
    end
    10'b 0101000001 : begin
      datar <= 16'b 0111010111110011;
      datai <= 16'b 1100111001001011;
      //65
    end
    10'b 0101000010 : begin
      datar <= 16'b 0111010110100101;
      datai <= 16'b 1100110110010010;
      //66
    end
    10'b 0101000011 : begin
      datar <= 16'b 0111010101010101;
      datai <= 16'b 1100110011011010;
      //67
    end
    10'b 0101000100 : begin
      datar <= 16'b 0111010100000100;
      datai <= 16'b 1100110000100001;
      //68
    end
    10'b 0101000101 : begin
      datar <= 16'b 0111010010110010;
      datai <= 16'b 1100101101101010;
      //69
    end
    10'b 0101000110 : begin
      datar <= 16'b 0111010001011111;
      datai <= 16'b 1100101010110011;
      //70
    end
    10'b 0101000111 : begin
      datar <= 16'b 0111010000001010;
      datai <= 16'b 1100100111111100;
      //71
    end
    10'b 0101001000 : begin
      datar <= 16'b 0111001110110101;
      datai <= 16'b 1100100101000110;
      //72
    end
    10'b 0101001001 : begin
      datar <= 16'b 0111001101011110;
      datai <= 16'b 1100100010010001;
      //73
    end
    10'b 0101001010 : begin
      datar <= 16'b 0111001100000111;
      datai <= 16'b 1100011111011100;
      //74
    end
    10'b 0101001011 : begin
      datar <= 16'b 0111001010101110;
      datai <= 16'b 1100011100100111;
      //75
    end
    10'b 0101001100 : begin
      datar <= 16'b 0111001001010100;
      datai <= 16'b 1100011001110100;
      //76
    end
    10'b 0101001101 : begin
      datar <= 16'b 0111000111111001;
      datai <= 16'b 1100010111000000;
      //77
    end
    10'b 0101001110 : begin
      datar <= 16'b 0111000110011101;
      datai <= 16'b 1100010100001110;
      //78
    end
    10'b 0101001111 : begin
      datar <= 16'b 0111000101000000;
      datai <= 16'b 1100010001011011;
      //79
    end
    10'b 0101010000 : begin
      datar <= 16'b 0111000011100010;
      datai <= 16'b 1100001110101010;
      //80
    end
    10'b 0101010001 : begin
      datar <= 16'b 0111000010000011;
      datai <= 16'b 1100001011111001;
      //81
    end
    10'b 0101010010 : begin
      datar <= 16'b 0111000000100010;
      datai <= 16'b 1100001001001000;
      //82
    end
    10'b 0101010011 : begin
      datar <= 16'b 0110111111000001;
      datai <= 16'b 1100000110011000;
      //83
    end
    10'b 0101010100 : begin
      datar <= 16'b 0110111101011110;
      datai <= 16'b 1100000011101001;
      //84
    end
    10'b 0101010101 : begin
      datar <= 16'b 0110111011111011;
      datai <= 16'b 1100000000111011;
      //85
    end
    10'b 0101010110 : begin
      datar <= 16'b 0110111010010110;
      datai <= 16'b 1011111110001101;
      //86
    end
    10'b 0101010111 : begin
      datar <= 16'b 0110111000110000;
      datai <= 16'b 1011111011011111;
      //87
    end
    10'b 0101011000 : begin
      datar <= 16'b 0110110111001001;
      datai <= 16'b 1011111000110010;
      //88
    end
    10'b 0101011001 : begin
      datar <= 16'b 0110110101100001;
      datai <= 16'b 1011110110000110;
      //89
    end
    10'b 0101011010 : begin
      datar <= 16'b 0110110011111000;
      datai <= 16'b 1011110011011011;
      //90
    end
    10'b 0101011011 : begin
      datar <= 16'b 0110110010001110;
      datai <= 16'b 1011110000110000;
      //91
    end
    10'b 0101011100 : begin
      datar <= 16'b 0110110000100011;
      datai <= 16'b 1011101110000110;
      //92
    end
    10'b 0101011101 : begin
      datar <= 16'b 0110101110110111;
      datai <= 16'b 1011101011011100;
      //93
    end
    10'b 0101011110 : begin
      datar <= 16'b 0110101101001010;
      datai <= 16'b 1011101000110011;
      //94
    end
    10'b 0101011111 : begin
      datar <= 16'b 0110101011011100;
      datai <= 16'b 1011100110001011;
      //95
    end
    10'b 0101100000 : begin
      datar <= 16'b 0110101001101101;
      datai <= 16'b 1011100011100100;
      //96
    end
    10'b 0101100001 : begin
      datar <= 16'b 0110100111111101;
      datai <= 16'b 1011100000111101;
      //97
    end
    10'b 0101100010 : begin
      datar <= 16'b 0110100110001011;
      datai <= 16'b 1011011110010111;
      //98
    end
    10'b 0101100011 : begin
      datar <= 16'b 0110100100011001;
      datai <= 16'b 1011011011110001;
      //99
    end
    10'b 0101100100 : begin
      datar <= 16'b 0110100010100110;
      datai <= 16'b 1011011001001100;
      //100
    end
    10'b 0101100101 : begin
      datar <= 16'b 0110100000110010;
      datai <= 16'b 1011010110101000;
      //101
    end
    10'b 0101100110 : begin
      datar <= 16'b 0110011110111100;
      datai <= 16'b 1011010100000101;
      //102
    end
    10'b 0101100111 : begin
      datar <= 16'b 0110011101000110;
      datai <= 16'b 1011010001100011;
      //103
    end
    10'b 0101101000 : begin
      datar <= 16'b 0110011011001111;
      datai <= 16'b 1011001111000001;
      //104
    end
    10'b 0101101001 : begin
      datar <= 16'b 0110011001010110;
      datai <= 16'b 1011001100100000;
      //105
    end
    10'b 0101101010 : begin
      datar <= 16'b 0110010111011101;
      datai <= 16'b 1011001001111111;
      //106
    end
    10'b 0101101011 : begin
      datar <= 16'b 0110010101100011;
      datai <= 16'b 1011000111100000;
      //107
    end
    10'b 0101101100 : begin
      datar <= 16'b 0110010011101000;
      datai <= 16'b 1011000101000001;
      //108
    end
    10'b 0101101101 : begin
      datar <= 16'b 0110010001101100;
      datai <= 16'b 1011000010100011;
      //109
    end
    10'b 0101101110 : begin
      datar <= 16'b 0110001111101110;
      datai <= 16'b 1011000000000101;
      //110
    end
    10'b 0101101111 : begin
      datar <= 16'b 0110001101110000;
      datai <= 16'b 1010111101101001;
      //111
    end
    10'b 0101110000 : begin
      datar <= 16'b 0110001011110001;
      datai <= 16'b 1010111011001101;
      //112
    end
    10'b 0101110001 : begin
      datar <= 16'b 0110001001110001;
      datai <= 16'b 1010111000110010;
      //113
    end
    10'b 0101110010 : begin
      datar <= 16'b 0110000111110000;
      datai <= 16'b 1010110110011000;
      //114
    end
    10'b 0101110011 : begin
      datar <= 16'b 0110000101101110;
      datai <= 16'b 1010110011111110;
      //115
    end
    10'b 0101110100 : begin
      datar <= 16'b 0110000011101011;
      datai <= 16'b 1010110001100101;
      //116
    end
    10'b 0101110101 : begin
      datar <= 16'b 0110000001101000;
      datai <= 16'b 1010101111001110;
      //117
    end
    10'b 0101110110 : begin
      datar <= 16'b 0101111111100011;
      datai <= 16'b 1010101100110111;
      //118
    end
    10'b 0101110111 : begin
      datar <= 16'b 0101111101011101;
      datai <= 16'b 1010101010100000;
      //119
    end
    10'b 0101111000 : begin
      datar <= 16'b 0101111011010111;
      datai <= 16'b 1010101000001011;
      //120
    end
    10'b 0101111001 : begin
      datar <= 16'b 0101111001001111;
      datai <= 16'b 1010100101110110;
      //121
    end
    10'b 0101111010 : begin
      datar <= 16'b 0101110111000111;
      datai <= 16'b 1010100011100011;
      //122
    end
    10'b 0101111011 : begin
      datar <= 16'b 0101110100111110;
      datai <= 16'b 1010100001010000;
      //123
    end
    10'b 0101111100 : begin
      datar <= 16'b 0101110010110011;
      datai <= 16'b 1010011110111110;
      //124
    end
    10'b 0101111101 : begin
      datar <= 16'b 0101110000101000;
      datai <= 16'b 1010011100101101;
      //125
    end
    10'b 0101111110 : begin
      datar <= 16'b 0101101110011100;
      datai <= 16'b 1010011010011100;
      //126
    end
    10'b 0101111111 : begin
      datar <= 16'b 0101101100001111;
      datai <= 16'b 1010011000001101;
      //127
    end
    10'b 0110000000 : begin
      datar <= 16'b 0101101010000010;
      datai <= 16'b 1010010101111110;
      //128
    end
    10'b 0110000001 : begin
      datar <= 16'b 0101100111110011;
      datai <= 16'b 1010010011110001;
      //129
    end
    10'b 0110000010 : begin
      datar <= 16'b 0101100101100100;
      datai <= 16'b 1010010001100100;
      //130
    end
    10'b 0110000011 : begin
      datar <= 16'b 0101100011010011;
      datai <= 16'b 1010001111011000;
      //131
    end
    10'b 0110000100 : begin
      datar <= 16'b 0101100001000010;
      datai <= 16'b 1010001101001101;
      //132
    end
    10'b 0110000101 : begin
      datar <= 16'b 0101011110110000;
      datai <= 16'b 1010001011000010;
      //133
    end
    10'b 0110000110 : begin
      datar <= 16'b 0101011100011101;
      datai <= 16'b 1010001000111001;
      //134
    end
    10'b 0110000111 : begin
      datar <= 16'b 0101011010001010;
      datai <= 16'b 1010000110110001;
      //135
    end
    10'b 0110001000 : begin
      datar <= 16'b 0101010111110101;
      datai <= 16'b 1010000100101001;
      //136
    end
    10'b 0110001001 : begin
      datar <= 16'b 0101010101100000;
      datai <= 16'b 1010000010100011;
      //137
    end
    10'b 0110001010 : begin
      datar <= 16'b 0101010011001001;
      datai <= 16'b 1010000000011101;
      //138
    end
    10'b 0110001011 : begin
      datar <= 16'b 0101010000110010;
      datai <= 16'b 1001111110011000;
      //139
    end
    10'b 0110001100 : begin
      datar <= 16'b 0101001110011011;
      datai <= 16'b 1001111100010101;
      //140
    end
    10'b 0110001101 : begin
      datar <= 16'b 0101001100000010;
      datai <= 16'b 1001111010010010;
      //141
    end
    10'b 0110001110 : begin
      datar <= 16'b 0101001001101000;
      datai <= 16'b 1001111000010000;
      //142
    end
    10'b 0110001111 : begin
      datar <= 16'b 0101000111001110;
      datai <= 16'b 1001110110001111;
      //143
    end
    10'b 0110010000 : begin
      datar <= 16'b 0101000100110011;
      datai <= 16'b 1001110100001111;
      //144
    end
    10'b 0110010001 : begin
      datar <= 16'b 0101000010010111;
      datai <= 16'b 1001110010010000;
      //145
    end
    10'b 0110010010 : begin
      datar <= 16'b 0100111111111011;
      datai <= 16'b 1001110000010010;
      //146
    end
    10'b 0110010011 : begin
      datar <= 16'b 0100111101011101;
      datai <= 16'b 1001101110010100;
      //147
    end
    10'b 0110010100 : begin
      datar <= 16'b 0100111010111111;
      datai <= 16'b 1001101100011000;
      //148
    end
    10'b 0110010101 : begin
      datar <= 16'b 0100111000100000;
      datai <= 16'b 1001101010011101;
      //149
    end
    10'b 0110010110 : begin
      datar <= 16'b 0100110110000001;
      datai <= 16'b 1001101000100011;
      //150
    end
    10'b 0110010111 : begin
      datar <= 16'b 0100110011100000;
      datai <= 16'b 1001100110101010;
      //151
    end
    10'b 0110011000 : begin
      datar <= 16'b 0100110000111111;
      datai <= 16'b 1001100100110001;
      //152
    end
    10'b 0110011001 : begin
      datar <= 16'b 0100101110011101;
      datai <= 16'b 1001100010111010;
      //153
    end
    10'b 0110011010 : begin
      datar <= 16'b 0100101011111011;
      datai <= 16'b 1001100001000100;
      //154
    end
    10'b 0110011011 : begin
      datar <= 16'b 0100101001011000;
      datai <= 16'b 1001011111001110;
      //155
    end
    10'b 0110011100 : begin
      datar <= 16'b 0100100110110100;
      datai <= 16'b 1001011101011010;
      //156
    end
    10'b 0110011101 : begin
      datar <= 16'b 0100100100001111;
      datai <= 16'b 1001011011100111;
      //157
    end
    10'b 0110011110 : begin
      datar <= 16'b 0100100001101001;
      datai <= 16'b 1001011001110101;
      //158
    end
    10'b 0110011111 : begin
      datar <= 16'b 0100011111000011;
      datai <= 16'b 1001011000000011;
      //159
    end
    10'b 0110100000 : begin
      datar <= 16'b 0100011100011100;
      datai <= 16'b 1001010110010011;
      //160
    end
    10'b 0110100001 : begin
      datar <= 16'b 0100011001110101;
      datai <= 16'b 1001010100100100;
      //161
    end
    10'b 0110100010 : begin
      datar <= 16'b 0100010111001101;
      datai <= 16'b 1001010010110110;
      //162
    end
    10'b 0110100011 : begin
      datar <= 16'b 0100010100100100;
      datai <= 16'b 1001010001001001;
      //163
    end
    10'b 0110100100 : begin
      datar <= 16'b 0100010001111010;
      datai <= 16'b 1001001111011101;
      //164
    end
    10'b 0110100101 : begin
      datar <= 16'b 0100001111010000;
      datai <= 16'b 1001001101110010;
      //165
    end
    10'b 0110100110 : begin
      datar <= 16'b 0100001100100101;
      datai <= 16'b 1001001100001000;
      //166
    end
    10'b 0110100111 : begin
      datar <= 16'b 0100001001111010;
      datai <= 16'b 1001001010011111;
      //167
    end
    10'b 0110101000 : begin
      datar <= 16'b 0100000111001110;
      datai <= 16'b 1001001000110111;
      //168
    end
    10'b 0110101001 : begin
      datar <= 16'b 0100000100100001;
      datai <= 16'b 1001000111010000;
      //169
    end
    10'b 0110101010 : begin
      datar <= 16'b 0100000001110011;
      datai <= 16'b 1001000101101010;
      //170
    end
    10'b 0110101011 : begin
      datar <= 16'b 0011111111000101;
      datai <= 16'b 1001000100000101;
      //171
    end
    10'b 0110101100 : begin
      datar <= 16'b 0011111100010111;
      datai <= 16'b 1001000010100010;
      //172
    end
    10'b 0110101101 : begin
      datar <= 16'b 0011111001101000;
      datai <= 16'b 1001000000111111;
      //173
    end
    10'b 0110101110 : begin
      datar <= 16'b 0011110110111000;
      datai <= 16'b 1000111111011110;
      //174
    end
    10'b 0110101111 : begin
      datar <= 16'b 0011110100000111;
      datai <= 16'b 1000111101111101;
      //175
    end
    10'b 0110110000 : begin
      datar <= 16'b 0011110001010110;
      datai <= 16'b 1000111100011110;
      //176
    end
    10'b 0110110001 : begin
      datar <= 16'b 0011101110100101;
      datai <= 16'b 1000111011000000;
      //177
    end
    10'b 0110110010 : begin
      datar <= 16'b 0011101011110010;
      datai <= 16'b 1000111001100011;
      //178
    end
    10'b 0110110011 : begin
      datar <= 16'b 0011101001000000;
      datai <= 16'b 1000111000000111;
      //179
    end
    10'b 0110110100 : begin
      datar <= 16'b 0011100110001100;
      datai <= 16'b 1000110110101100;
      //180
    end
    10'b 0110110101 : begin
      datar <= 16'b 0011100011011001;
      datai <= 16'b 1000110101010010;
      //181
    end
    10'b 0110110110 : begin
      datar <= 16'b 0011100000100100;
      datai <= 16'b 1000110011111001;
      //182
    end
    10'b 0110110111 : begin
      datar <= 16'b 0011011101101111;
      datai <= 16'b 1000110010100010;
      //183
    end
    10'b 0110111000 : begin
      datar <= 16'b 0011011010111010;
      datai <= 16'b 1000110001001011;
      //184
    end
    10'b 0110111001 : begin
      datar <= 16'b 0011011000000100;
      datai <= 16'b 1000101111110110;
      //185
    end
    10'b 0110111010 : begin
      datar <= 16'b 0011010101001101;
      datai <= 16'b 1000101110100001;
      //186
    end
    10'b 0110111011 : begin
      datar <= 16'b 0011010010010110;
      datai <= 16'b 1000101101001110;
      //187
    end
    10'b 0110111100 : begin
      datar <= 16'b 0011001111011111;
      datai <= 16'b 1000101011111100;
      //188
    end
    10'b 0110111101 : begin
      datar <= 16'b 0011001100100110;
      datai <= 16'b 1000101010101011;
      //189
    end
    10'b 0110111110 : begin
      datar <= 16'b 0011001001101110;
      datai <= 16'b 1000101001011011;
      //190
    end
    10'b 0110111111 : begin
      datar <= 16'b 0011000110110101;
      datai <= 16'b 1000101000001101;
      //191
    end
    10'b 0111000000 : begin
      datar <= 16'b 0011000011111011;
      datai <= 16'b 1000100110111111;
      //192
    end
    10'b 0111000001 : begin
      datar <= 16'b 0011000001000001;
      datai <= 16'b 1000100101110011;
      //193
    end
    10'b 0111000010 : begin
      datar <= 16'b 0010111110000111;
      datai <= 16'b 1000100100101000;
      //194
    end
    10'b 0111000011 : begin
      datar <= 16'b 0010111011001100;
      datai <= 16'b 1000100011011110;
      //195
    end
    10'b 0111000100 : begin
      datar <= 16'b 0010111000010001;
      datai <= 16'b 1000100010010101;
      //196
    end
    10'b 0111000101 : begin
      datar <= 16'b 0010110101010101;
      datai <= 16'b 1000100001001101;
      //197
    end
    10'b 0111000110 : begin
      datar <= 16'b 0010110010011001;
      datai <= 16'b 1000100000000110;
      //198
    end
    10'b 0111000111 : begin
      datar <= 16'b 0010101111011100;
      datai <= 16'b 1000011111000001;
      //199
    end
    10'b 0111001000 : begin
      datar <= 16'b 0010101100011111;
      datai <= 16'b 1000011101111100;
      //200
    end
    10'b 0111001001 : begin
      datar <= 16'b 0010101001100001;
      datai <= 16'b 1000011100111001;
      //201
    end
    10'b 0111001010 : begin
      datar <= 16'b 0010100110100011;
      datai <= 16'b 1000011011110111;
      //202
    end
    10'b 0111001011 : begin
      datar <= 16'b 0010100011100101;
      datai <= 16'b 1000011010110110;
      //203
    end
    10'b 0111001100 : begin
      datar <= 16'b 0010100000100110;
      datai <= 16'b 1000011001110111;
      //204
    end
    10'b 0111001101 : begin
      datar <= 16'b 0010011101100111;
      datai <= 16'b 1000011000111000;
      //205
    end
    10'b 0111001110 : begin
      datar <= 16'b 0010011010101000;
      datai <= 16'b 1000010111111011;
      //206
    end
    10'b 0111001111 : begin
      datar <= 16'b 0010010111101000;
      datai <= 16'b 1000010110111111;
      //207
    end
    10'b 0111010000 : begin
      datar <= 16'b 0010010100101000;
      datai <= 16'b 1000010110000100;
      //208
    end
    10'b 0111010001 : begin
      datar <= 16'b 0010010001100111;
      datai <= 16'b 1000010101001010;
      //209
    end
    10'b 0111010010 : begin
      datar <= 16'b 0010001110100110;
      datai <= 16'b 1000010100010010;
      //210
    end
    10'b 0111010011 : begin
      datar <= 16'b 0010001011100101;
      datai <= 16'b 1000010011011010;
      //211
    end
    10'b 0111010100 : begin
      datar <= 16'b 0010001000100011;
      datai <= 16'b 1000010010100100;
      //212
    end
    10'b 0111010101 : begin
      datar <= 16'b 0010000101100001;
      datai <= 16'b 1000010001101111;
      //213
    end
    10'b 0111010110 : begin
      datar <= 16'b 0010000010011111;
      datai <= 16'b 1000010000111011;
      //214
    end
    10'b 0111010111 : begin
      datar <= 16'b 0001111111011101;
      datai <= 16'b 1000010000001000;
      //215
    end
    10'b 0111011000 : begin
      datar <= 16'b 0001111100011010;
      datai <= 16'b 1000001111010111;
      //216
    end
    10'b 0111011001 : begin
      datar <= 16'b 0001111001010111;
      datai <= 16'b 1000001110100111;
      //217
    end
    10'b 0111011010 : begin
      datar <= 16'b 0001110110010011;
      datai <= 16'b 1000001101111000;
      //218
    end
    10'b 0111011011 : begin
      datar <= 16'b 0001110011001111;
      datai <= 16'b 1000001101001010;
      //219
    end
    10'b 0111011100 : begin
      datar <= 16'b 0001110000001011;
      datai <= 16'b 1000001100011101;
      //220
    end
    10'b 0111011101 : begin
      datar <= 16'b 0001101101000111;
      datai <= 16'b 1000001011110010;
      //221
    end
    10'b 0111011110 : begin
      datar <= 16'b 0001101010000010;
      datai <= 16'b 1000001011000111;
      //222
    end
    10'b 0111011111 : begin
      datar <= 16'b 0001100110111110;
      datai <= 16'b 1000001010011110;
      //223
    end
    10'b 0111100000 : begin
      datar <= 16'b 0001100011111001;
      datai <= 16'b 1000001001110111;
      //224
    end
    10'b 0111100001 : begin
      datar <= 16'b 0001100000110011;
      datai <= 16'b 1000001001010000;
      //225
    end
    10'b 0111100010 : begin
      datar <= 16'b 0001011101101110;
      datai <= 16'b 1000001000101011;
      //226
    end
    10'b 0111100011 : begin
      datar <= 16'b 0001011010101000;
      datai <= 16'b 1000001000000110;
      //227
    end
    10'b 0111100100 : begin
      datar <= 16'b 0001010111100010;
      datai <= 16'b 1000000111100011;
      //228
    end
    10'b 0111100101 : begin
      datar <= 16'b 0001010100011100;
      datai <= 16'b 1000000111000010;
      //229
    end
    10'b 0111100110 : begin
      datar <= 16'b 0001010001010101;
      datai <= 16'b 1000000110100001;
      //230
    end
    10'b 0111100111 : begin
      datar <= 16'b 0001001110001111;
      datai <= 16'b 1000000110000010;
      //231
    end
    10'b 0111101000 : begin
      datar <= 16'b 0001001011001000;
      datai <= 16'b 1000000101100100;
      //232
    end
    10'b 0111101001 : begin
      datar <= 16'b 0001001000000001;
      datai <= 16'b 1000000101000111;
      //233
    end
    10'b 0111101010 : begin
      datar <= 16'b 0001000100111010;
      datai <= 16'b 1000000100101011;
      //234
    end
    10'b 0111101011 : begin
      datar <= 16'b 0001000001110010;
      datai <= 16'b 1000000100010001;
      //235
    end
    10'b 0111101100 : begin
      datar <= 16'b 0000111110101011;
      datai <= 16'b 1000000011110111;
      //236
    end
    10'b 0111101101 : begin
      datar <= 16'b 0000111011100011;
      datai <= 16'b 1000000011011111;
      //237
    end
    10'b 0111101110 : begin
      datar <= 16'b 0000111000011100;
      datai <= 16'b 1000000011001001;
      //238
    end
    10'b 0111101111 : begin
      datar <= 16'b 0000110101010100;
      datai <= 16'b 1000000010110011;
      //239
    end
    10'b 0111110000 : begin
      datar <= 16'b 0000110010001100;
      datai <= 16'b 1000000010011111;
      //240
    end
    10'b 0111110001 : begin
      datar <= 16'b 0000101111000100;
      datai <= 16'b 1000000010001100;
      //241
    end
    10'b 0111110010 : begin
      datar <= 16'b 0000101011111011;
      datai <= 16'b 1000000001111010;
      //242
    end
    10'b 0111110011 : begin
      datar <= 16'b 0000101000110011;
      datai <= 16'b 1000000001101001;
      //243
    end
    10'b 0111110100 : begin
      datar <= 16'b 0000100101101010;
      datai <= 16'b 1000000001011010;
      //244
    end
    10'b 0111110101 : begin
      datar <= 16'b 0000100010100010;
      datai <= 16'b 1000000001001100;
      //245
    end
    10'b 0111110110 : begin
      datar <= 16'b 0000011111011001;
      datai <= 16'b 1000000000111111;
      //246
    end
    10'b 0111110111 : begin
      datar <= 16'b 0000011100010001;
      datai <= 16'b 1000000000110011;
      //247
    end
    10'b 0111111000 : begin
      datar <= 16'b 0000011001001000;
      datai <= 16'b 1000000000101000;
      //248
    end
    10'b 0111111001 : begin
      datar <= 16'b 0000010101111111;
      datai <= 16'b 1000000000011111;
      //249
    end
    10'b 0111111010 : begin
      datar <= 16'b 0000010010110110;
      datai <= 16'b 1000000000010111;
      //250
    end
    10'b 0111111011 : begin
      datar <= 16'b 0000001111101101;
      datai <= 16'b 1000000000010000;
      //251
    end
    10'b 0111111100 : begin
      datar <= 16'b 0000001100100100;
      datai <= 16'b 1000000000001011;
      //252
    end
    10'b 0111111101 : begin
      datar <= 16'b 0000001001011011;
      datai <= 16'b 1000000000000111;
      //253
    end
    10'b 0111111110 : begin
      datar <= 16'b 0000000110010010;
      datai <= 16'b 1000000000000011;
      //254
    end
    10'b 0111111111 : begin
      datar <= 16'b 0000000011001001;
      datai <= 16'b 1000000000000010;
      //255
    end
    10'b 1000000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1000000001 : begin
      datar <= 16'b 0111111111111001;
      datai <= 16'b 1111110110100101;
      //3
    end
    10'b 1000000010 : begin
      datar <= 16'b 0111111111101001;
      datai <= 16'b 1111101101001010;
      //6
    end
    10'b 1000000011 : begin
      datar <= 16'b 0111111111001101;
      datai <= 16'b 1111100011101111;
      //9
    end
    10'b 1000000100 : begin
      datar <= 16'b 0111111110100110;
      datai <= 16'b 1111011010010110;
      //12
    end
    10'b 1000000101 : begin
      datar <= 16'b 0111111101110100;
      datai <= 16'b 1111010000111100;
      //15
    end
    10'b 1000000110 : begin
      datar <= 16'b 0111111100110111;
      datai <= 16'b 1111000111100100;
      //18
    end
    10'b 1000000111 : begin
      datar <= 16'b 0111111011101111;
      datai <= 16'b 1110111110001110;
      //21
    end
    10'b 1000001000 : begin
      datar <= 16'b 0111111010011100;
      datai <= 16'b 1110110100111000;
      //24
    end
    10'b 1000001001 : begin
      datar <= 16'b 0111111000111110;
      datai <= 16'b 1110101011100100;
      //27
    end
    10'b 1000001010 : begin
      datar <= 16'b 0111110111010101;
      datai <= 16'b 1110100010010010;
      //30
    end
    10'b 1000001011 : begin
      datar <= 16'b 0111110101100010;
      datai <= 16'b 1110011001000010;
      //33
    end
    10'b 1000001100 : begin
      datar <= 16'b 0111110011100011;
      datai <= 16'b 1110001111110101;
      //36
    end
    10'b 1000001101 : begin
      datar <= 16'b 0111110001011001;
      datai <= 16'b 1110000110101001;
      //39
    end
    10'b 1000001110 : begin
      datar <= 16'b 0111101111000101;
      datai <= 16'b 1101111101100001;
      //42
    end
    10'b 1000001111 : begin
      datar <= 16'b 0111101100100110;
      datai <= 16'b 1101110100011011;
      //45
    end
    10'b 1000010000 : begin
      datar <= 16'b 0111101001111100;
      datai <= 16'b 1101101011011000;
      //48
    end
    10'b 1000010001 : begin
      datar <= 16'b 0111100111001000;
      datai <= 16'b 1101100010011001;
      //51
    end
    10'b 1000010010 : begin
      datar <= 16'b 0111100100001001;
      datai <= 16'b 1101011001011101;
      //54
    end
    10'b 1000010011 : begin
      datar <= 16'b 0111100000111111;
      datai <= 16'b 1101010000100100;
      //57
    end
    10'b 1000010100 : begin
      datar <= 16'b 0111011101101011;
      datai <= 16'b 1101000111101111;
      //60
    end
    10'b 1000010101 : begin
      datar <= 16'b 0111011010001101;
      datai <= 16'b 1100111110111111;
      //63
    end
    10'b 1000010110 : begin
      datar <= 16'b 0111010110100101;
      datai <= 16'b 1100110110010010;
      //66
    end
    10'b 1000010111 : begin
      datar <= 16'b 0111010010110010;
      datai <= 16'b 1100101101101010;
      //69
    end
    10'b 1000011000 : begin
      datar <= 16'b 0111001110110101;
      datai <= 16'b 1100100101000110;
      //72
    end
    10'b 1000011001 : begin
      datar <= 16'b 0111001010101110;
      datai <= 16'b 1100011100100111;
      //75
    end
    10'b 1000011010 : begin
      datar <= 16'b 0111000110011101;
      datai <= 16'b 1100010100001110;
      //78
    end
    10'b 1000011011 : begin
      datar <= 16'b 0111000010000011;
      datai <= 16'b 1100001011111001;
      //81
    end
    10'b 1000011100 : begin
      datar <= 16'b 0110111101011110;
      datai <= 16'b 1100000011101001;
      //84
    end
    10'b 1000011101 : begin
      datar <= 16'b 0110111000110000;
      datai <= 16'b 1011111011011111;
      //87
    end
    10'b 1000011110 : begin
      datar <= 16'b 0110110011111000;
      datai <= 16'b 1011110011011011;
      //90
    end
    10'b 1000011111 : begin
      datar <= 16'b 0110101110110111;
      datai <= 16'b 1011101011011100;
      //93
    end
    10'b 1000100000 : begin
      datar <= 16'b 0110101001101101;
      datai <= 16'b 1011100011100100;
      //96
    end
    10'b 1000100001 : begin
      datar <= 16'b 0110100100011001;
      datai <= 16'b 1011011011110001;
      //99
    end
    10'b 1000100010 : begin
      datar <= 16'b 0110011110111100;
      datai <= 16'b 1011010100000101;
      //102
    end
    10'b 1000100011 : begin
      datar <= 16'b 0110011001010110;
      datai <= 16'b 1011001100100000;
      //105
    end
    10'b 1000100100 : begin
      datar <= 16'b 0110010011101000;
      datai <= 16'b 1011000101000001;
      //108
    end
    10'b 1000100101 : begin
      datar <= 16'b 0110001101110000;
      datai <= 16'b 1010111101101001;
      //111
    end
    10'b 1000100110 : begin
      datar <= 16'b 0110000111110000;
      datai <= 16'b 1010110110011000;
      //114
    end
    10'b 1000100111 : begin
      datar <= 16'b 0110000001101000;
      datai <= 16'b 1010101111001110;
      //117
    end
    10'b 1000101000 : begin
      datar <= 16'b 0101111011010111;
      datai <= 16'b 1010101000001011;
      //120
    end
    10'b 1000101001 : begin
      datar <= 16'b 0101110100111110;
      datai <= 16'b 1010100001010000;
      //123
    end
    10'b 1000101010 : begin
      datar <= 16'b 0101101110011100;
      datai <= 16'b 1010011010011100;
      //126
    end
    10'b 1000101011 : begin
      datar <= 16'b 0101100111110011;
      datai <= 16'b 1010010011110001;
      //129
    end
    10'b 1000101100 : begin
      datar <= 16'b 0101100001000010;
      datai <= 16'b 1010001101001101;
      //132
    end
    10'b 1000101101 : begin
      datar <= 16'b 0101011010001010;
      datai <= 16'b 1010000110110001;
      //135
    end
    10'b 1000101110 : begin
      datar <= 16'b 0101010011001001;
      datai <= 16'b 1010000000011101;
      //138
    end
    10'b 1000101111 : begin
      datar <= 16'b 0101001100000010;
      datai <= 16'b 1001111010010010;
      //141
    end
    10'b 1000110000 : begin
      datar <= 16'b 0101000100110011;
      datai <= 16'b 1001110100001111;
      //144
    end
    10'b 1000110001 : begin
      datar <= 16'b 0100111101011101;
      datai <= 16'b 1001101110010100;
      //147
    end
    10'b 1000110010 : begin
      datar <= 16'b 0100110110000001;
      datai <= 16'b 1001101000100011;
      //150
    end
    10'b 1000110011 : begin
      datar <= 16'b 0100101110011101;
      datai <= 16'b 1001100010111010;
      //153
    end
    10'b 1000110100 : begin
      datar <= 16'b 0100100110110100;
      datai <= 16'b 1001011101011010;
      //156
    end
    10'b 1000110101 : begin
      datar <= 16'b 0100011111000011;
      datai <= 16'b 1001011000000011;
      //159
    end
    10'b 1000110110 : begin
      datar <= 16'b 0100010111001101;
      datai <= 16'b 1001010010110110;
      //162
    end
    10'b 1000110111 : begin
      datar <= 16'b 0100001111010000;
      datai <= 16'b 1001001101110010;
      //165
    end
    10'b 1000111000 : begin
      datar <= 16'b 0100000111001110;
      datai <= 16'b 1001001000110111;
      //168
    end
    10'b 1000111001 : begin
      datar <= 16'b 0011111111000101;
      datai <= 16'b 1001000100000101;
      //171
    end
    10'b 1000111010 : begin
      datar <= 16'b 0011110110111000;
      datai <= 16'b 1000111111011110;
      //174
    end
    10'b 1000111011 : begin
      datar <= 16'b 0011101110100101;
      datai <= 16'b 1000111011000000;
      //177
    end
    10'b 1000111100 : begin
      datar <= 16'b 0011100110001100;
      datai <= 16'b 1000110110101100;
      //180
    end
    10'b 1000111101 : begin
      datar <= 16'b 0011011101101111;
      datai <= 16'b 1000110010100010;
      //183
    end
    10'b 1000111110 : begin
      datar <= 16'b 0011010101001101;
      datai <= 16'b 1000101110100001;
      //186
    end
    10'b 1000111111 : begin
      datar <= 16'b 0011001100100110;
      datai <= 16'b 1000101010101011;
      //189
    end
    10'b 1001000000 : begin
      datar <= 16'b 0011000011111011;
      datai <= 16'b 1000100110111111;
      //192
    end
    10'b 1001000001 : begin
      datar <= 16'b 0010111011001100;
      datai <= 16'b 1000100011011110;
      //195
    end
    10'b 1001000010 : begin
      datar <= 16'b 0010110010011001;
      datai <= 16'b 1000100000000110;
      //198
    end
    10'b 1001000011 : begin
      datar <= 16'b 0010101001100001;
      datai <= 16'b 1000011100111001;
      //201
    end
    10'b 1001000100 : begin
      datar <= 16'b 0010100000100110;
      datai <= 16'b 1000011001110111;
      //204
    end
    10'b 1001000101 : begin
      datar <= 16'b 0010010111101000;
      datai <= 16'b 1000010110111111;
      //207
    end
    10'b 1001000110 : begin
      datar <= 16'b 0010001110100110;
      datai <= 16'b 1000010100010010;
      //210
    end
    10'b 1001000111 : begin
      datar <= 16'b 0010000101100001;
      datai <= 16'b 1000010001101111;
      //213
    end
    10'b 1001001000 : begin
      datar <= 16'b 0001111100011010;
      datai <= 16'b 1000001111010111;
      //216
    end
    10'b 1001001001 : begin
      datar <= 16'b 0001110011001111;
      datai <= 16'b 1000001101001010;
      //219
    end
    10'b 1001001010 : begin
      datar <= 16'b 0001101010000010;
      datai <= 16'b 1000001011000111;
      //222
    end
    10'b 1001001011 : begin
      datar <= 16'b 0001100000110011;
      datai <= 16'b 1000001001010000;
      //225
    end
    10'b 1001001100 : begin
      datar <= 16'b 0001010111100010;
      datai <= 16'b 1000000111100011;
      //228
    end
    10'b 1001001101 : begin
      datar <= 16'b 0001001110001111;
      datai <= 16'b 1000000110000010;
      //231
    end
    10'b 1001001110 : begin
      datar <= 16'b 0001000100111010;
      datai <= 16'b 1000000100101011;
      //234
    end
    10'b 1001001111 : begin
      datar <= 16'b 0000111011100011;
      datai <= 16'b 1000000011011111;
      //237
    end
    10'b 1001010000 : begin
      datar <= 16'b 0000110010001100;
      datai <= 16'b 1000000010011111;
      //240
    end
    10'b 1001010001 : begin
      datar <= 16'b 0000101000110011;
      datai <= 16'b 1000000001101001;
      //243
    end
    10'b 1001010010 : begin
      datar <= 16'b 0000011111011001;
      datai <= 16'b 1000000000111111;
      //246
    end
    10'b 1001010011 : begin
      datar <= 16'b 0000010101111111;
      datai <= 16'b 1000000000011111;
      //249
    end
    10'b 1001010100 : begin
      datar <= 16'b 0000001100100100;
      datai <= 16'b 1000000000001011;
      //252
    end
    10'b 1001010101 : begin
      datar <= 16'b 0000000011001001;
      datai <= 16'b 1000000000000010;
      //255
    end
    10'b 1001010110 : begin
      datar <= 16'b 1111111001101110;
      datai <= 16'b 1000000000000011;
      //258
    end
    10'b 1001010111 : begin
      datar <= 16'b 1111110000010011;
      datai <= 16'b 1000000000010000;
      //261
    end
    10'b 1001011000 : begin
      datar <= 16'b 1111100110111000;
      datai <= 16'b 1000000000101000;
      //264
    end
    10'b 1001011001 : begin
      datar <= 16'b 1111011101011110;
      datai <= 16'b 1000000001001100;
      //267
    end
    10'b 1001011010 : begin
      datar <= 16'b 1111010100000101;
      datai <= 16'b 1000000001111010;
      //270
    end
    10'b 1001011011 : begin
      datar <= 16'b 1111001010101100;
      datai <= 16'b 1000000010110011;
      //273
    end
    10'b 1001011100 : begin
      datar <= 16'b 1111000001010101;
      datai <= 16'b 1000000011110111;
      //276
    end
    10'b 1001011101 : begin
      datar <= 16'b 1110110111111111;
      datai <= 16'b 1000000101000111;
      //279
    end
    10'b 1001011110 : begin
      datar <= 16'b 1110101110101011;
      datai <= 16'b 1000000110100001;
      //282
    end
    10'b 1001011111 : begin
      datar <= 16'b 1110100101011000;
      datai <= 16'b 1000001000000110;
      //285
    end
    10'b 1001100000 : begin
      datar <= 16'b 1110011100000111;
      datai <= 16'b 1000001001110111;
      //288
    end
    10'b 1001100001 : begin
      datar <= 16'b 1110010010111001;
      datai <= 16'b 1000001011110010;
      //291
    end
    10'b 1001100010 : begin
      datar <= 16'b 1110001001101101;
      datai <= 16'b 1000001101111000;
      //294
    end
    10'b 1001100011 : begin
      datar <= 16'b 1110000000100011;
      datai <= 16'b 1000010000001000;
      //297
    end
    10'b 1001100100 : begin
      datar <= 16'b 1101110111011101;
      datai <= 16'b 1000010010100100;
      //300
    end
    10'b 1001100101 : begin
      datar <= 16'b 1101101110011001;
      datai <= 16'b 1000010101001010;
      //303
    end
    10'b 1001100110 : begin
      datar <= 16'b 1101100101011000;
      datai <= 16'b 1000010111111011;
      //306
    end
    10'b 1001100111 : begin
      datar <= 16'b 1101011100011011;
      datai <= 16'b 1000011010110110;
      //309
    end
    10'b 1001101000 : begin
      datar <= 16'b 1101010011100001;
      datai <= 16'b 1000011101111100;
      //312
    end
    10'b 1001101001 : begin
      datar <= 16'b 1101001010101011;
      datai <= 16'b 1000100001001101;
      //315
    end
    10'b 1001101010 : begin
      datar <= 16'b 1101000001111001;
      datai <= 16'b 1000100100101000;
      //318
    end
    10'b 1001101011 : begin
      datar <= 16'b 1100111001001011;
      datai <= 16'b 1000101000001101;
      //321
    end
    10'b 1001101100 : begin
      datar <= 16'b 1100110000100001;
      datai <= 16'b 1000101011111100;
      //324
    end
    10'b 1001101101 : begin
      datar <= 16'b 1100100111111100;
      datai <= 16'b 1000101111110110;
      //327
    end
    10'b 1001101110 : begin
      datar <= 16'b 1100011111011100;
      datai <= 16'b 1000110011111001;
      //330
    end
    10'b 1001101111 : begin
      datar <= 16'b 1100010111000000;
      datai <= 16'b 1000111000000111;
      //333
    end
    10'b 1001110000 : begin
      datar <= 16'b 1100001110101010;
      datai <= 16'b 1000111100011110;
      //336
    end
    10'b 1001110001 : begin
      datar <= 16'b 1100000110011000;
      datai <= 16'b 1001000000111111;
      //339
    end
    10'b 1001110010 : begin
      datar <= 16'b 1011111110001101;
      datai <= 16'b 1001000101101010;
      //342
    end
    10'b 1001110011 : begin
      datar <= 16'b 1011110110000110;
      datai <= 16'b 1001001010011111;
      //345
    end
    10'b 1001110100 : begin
      datar <= 16'b 1011101110000110;
      datai <= 16'b 1001001111011101;
      //348
    end
    10'b 1001110101 : begin
      datar <= 16'b 1011100110001011;
      datai <= 16'b 1001010100100100;
      //351
    end
    10'b 1001110110 : begin
      datar <= 16'b 1011011110010111;
      datai <= 16'b 1001011001110101;
      //354
    end
    10'b 1001110111 : begin
      datar <= 16'b 1011010110101000;
      datai <= 16'b 1001011111001110;
      //357
    end
    10'b 1001111000 : begin
      datar <= 16'b 1011001111000001;
      datai <= 16'b 1001100100110001;
      //360
    end
    10'b 1001111001 : begin
      datar <= 16'b 1011000111100000;
      datai <= 16'b 1001101010011101;
      //363
    end
    10'b 1001111010 : begin
      datar <= 16'b 1011000000000101;
      datai <= 16'b 1001110000010010;
      //366
    end
    10'b 1001111011 : begin
      datar <= 16'b 1010111000110010;
      datai <= 16'b 1001110110001111;
      //369
    end
    10'b 1001111100 : begin
      datar <= 16'b 1010110001100101;
      datai <= 16'b 1001111100010101;
      //372
    end
    10'b 1001111101 : begin
      datar <= 16'b 1010101010100000;
      datai <= 16'b 1010000010100011;
      //375
    end
    10'b 1001111110 : begin
      datar <= 16'b 1010100011100011;
      datai <= 16'b 1010001000111001;
      //378
    end
    10'b 1001111111 : begin
      datar <= 16'b 1010011100101101;
      datai <= 16'b 1010001111011000;
      //381
    end
    10'b 1010000000 : begin
      datar <= 16'b 1010010101111110;
      datai <= 16'b 1010010101111110;
      //384
    end
    10'b 1010000001 : begin
      datar <= 16'b 1010001111011000;
      datai <= 16'b 1010011100101101;
      //387
    end
    10'b 1010000010 : begin
      datar <= 16'b 1010001000111001;
      datai <= 16'b 1010100011100011;
      //390
    end
    10'b 1010000011 : begin
      datar <= 16'b 1010000010100011;
      datai <= 16'b 1010101010100000;
      //393
    end
    10'b 1010000100 : begin
      datar <= 16'b 1001111100010101;
      datai <= 16'b 1010110001100101;
      //396
    end
    10'b 1010000101 : begin
      datar <= 16'b 1001110110001111;
      datai <= 16'b 1010111000110010;
      //399
    end
    10'b 1010000110 : begin
      datar <= 16'b 1001110000010010;
      datai <= 16'b 1011000000000101;
      //402
    end
    10'b 1010000111 : begin
      datar <= 16'b 1001101010011101;
      datai <= 16'b 1011000111100000;
      //405
    end
    10'b 1010001000 : begin
      datar <= 16'b 1001100100110001;
      datai <= 16'b 1011001111000001;
      //408
    end
    10'b 1010001001 : begin
      datar <= 16'b 1001011111001110;
      datai <= 16'b 1011010110101000;
      //411
    end
    10'b 1010001010 : begin
      datar <= 16'b 1001011001110101;
      datai <= 16'b 1011011110010111;
      //414
    end
    10'b 1010001011 : begin
      datar <= 16'b 1001010100100100;
      datai <= 16'b 1011100110001011;
      //417
    end
    10'b 1010001100 : begin
      datar <= 16'b 1001001111011101;
      datai <= 16'b 1011101110000110;
      //420
    end
    10'b 1010001101 : begin
      datar <= 16'b 1001001010011111;
      datai <= 16'b 1011110110000110;
      //423
    end
    10'b 1010001110 : begin
      datar <= 16'b 1001000101101010;
      datai <= 16'b 1011111110001101;
      //426
    end
    10'b 1010001111 : begin
      datar <= 16'b 1001000000111111;
      datai <= 16'b 1100000110011000;
      //429
    end
    10'b 1010010000 : begin
      datar <= 16'b 1000111100011110;
      datai <= 16'b 1100001110101010;
      //432
    end
    10'b 1010010001 : begin
      datar <= 16'b 1000111000000111;
      datai <= 16'b 1100010111000000;
      //435
    end
    10'b 1010010010 : begin
      datar <= 16'b 1000110011111001;
      datai <= 16'b 1100011111011100;
      //438
    end
    10'b 1010010011 : begin
      datar <= 16'b 1000101111110110;
      datai <= 16'b 1100100111111100;
      //441
    end
    10'b 1010010100 : begin
      datar <= 16'b 1000101011111100;
      datai <= 16'b 1100110000100001;
      //444
    end
    10'b 1010010101 : begin
      datar <= 16'b 1000101000001101;
      datai <= 16'b 1100111001001011;
      //447
    end
    10'b 1010010110 : begin
      datar <= 16'b 1000100100101000;
      datai <= 16'b 1101000001111001;
      //450
    end
    10'b 1010010111 : begin
      datar <= 16'b 1000100001001101;
      datai <= 16'b 1101001010101011;
      //453
    end
    10'b 1010011000 : begin
      datar <= 16'b 1000011101111100;
      datai <= 16'b 1101010011100001;
      //456
    end
    10'b 1010011001 : begin
      datar <= 16'b 1000011010110110;
      datai <= 16'b 1101011100011011;
      //459
    end
    10'b 1010011010 : begin
      datar <= 16'b 1000010111111011;
      datai <= 16'b 1101100101011000;
      //462
    end
    10'b 1010011011 : begin
      datar <= 16'b 1000010101001010;
      datai <= 16'b 1101101110011001;
      //465
    end
    10'b 1010011100 : begin
      datar <= 16'b 1000010010100100;
      datai <= 16'b 1101110111011101;
      //468
    end
    10'b 1010011101 : begin
      datar <= 16'b 1000010000001000;
      datai <= 16'b 1110000000100011;
      //471
    end
    10'b 1010011110 : begin
      datar <= 16'b 1000001101111000;
      datai <= 16'b 1110001001101101;
      //474
    end
    10'b 1010011111 : begin
      datar <= 16'b 1000001011110010;
      datai <= 16'b 1110010010111001;
      //477
    end
    10'b 1010100000 : begin
      datar <= 16'b 1000001001110111;
      datai <= 16'b 1110011100000111;
      //480
    end
    10'b 1010100001 : begin
      datar <= 16'b 1000001000000110;
      datai <= 16'b 1110100101011000;
      //483
    end
    10'b 1010100010 : begin
      datar <= 16'b 1000000110100001;
      datai <= 16'b 1110101110101011;
      //486
    end
    10'b 1010100011 : begin
      datar <= 16'b 1000000101000111;
      datai <= 16'b 1110110111111111;
      //489
    end
    10'b 1010100100 : begin
      datar <= 16'b 1000000011110111;
      datai <= 16'b 1111000001010101;
      //492
    end
    10'b 1010100101 : begin
      datar <= 16'b 1000000010110011;
      datai <= 16'b 1111001010101100;
      //495
    end
    10'b 1010100110 : begin
      datar <= 16'b 1000000001111010;
      datai <= 16'b 1111010100000101;
      //498
    end
    10'b 1010100111 : begin
      datar <= 16'b 1000000001001100;
      datai <= 16'b 1111011101011110;
      //501
    end
    10'b 1010101000 : begin
      datar <= 16'b 1000000000101000;
      datai <= 16'b 1111100110111000;
      //504
    end
    10'b 1010101001 : begin
      datar <= 16'b 1000000000010000;
      datai <= 16'b 1111110000010011;
      //507
    end
    10'b 1010101010 : begin
      datar <= 16'b 1000000000000011;
      datai <= 16'b 1111111001101110;
      //510
    end
    10'b 1010101011 : begin
      datar <= 16'b 1000000000000010;
      datai <= 16'b 0000000011001001;
      //513
    end
    10'b 1010101100 : begin
      datar <= 16'b 1000000000001011;
      datai <= 16'b 0000001100100100;
      //516
    end
    10'b 1010101101 : begin
      datar <= 16'b 1000000000011111;
      datai <= 16'b 0000010101111111;
      //519
    end
    10'b 1010101110 : begin
      datar <= 16'b 1000000000111111;
      datai <= 16'b 0000011111011001;
      //522
    end
    10'b 1010101111 : begin
      datar <= 16'b 1000000001101001;
      datai <= 16'b 0000101000110011;
      //525
    end
    10'b 1010110000 : begin
      datar <= 16'b 1000000010011111;
      datai <= 16'b 0000110010001100;
      //528
    end
    10'b 1010110001 : begin
      datar <= 16'b 1000000011011111;
      datai <= 16'b 0000111011100011;
      //531
    end
    10'b 1010110010 : begin
      datar <= 16'b 1000000100101011;
      datai <= 16'b 0001000100111010;
      //534
    end
    10'b 1010110011 : begin
      datar <= 16'b 1000000110000010;
      datai <= 16'b 0001001110001111;
      //537
    end
    10'b 1010110100 : begin
      datar <= 16'b 1000000111100011;
      datai <= 16'b 0001010111100010;
      //540
    end
    10'b 1010110101 : begin
      datar <= 16'b 1000001001010000;
      datai <= 16'b 0001100000110011;
      //543
    end
    10'b 1010110110 : begin
      datar <= 16'b 1000001011000111;
      datai <= 16'b 0001101010000010;
      //546
    end
    10'b 1010110111 : begin
      datar <= 16'b 1000001101001010;
      datai <= 16'b 0001110011001111;
      //549
    end
    10'b 1010111000 : begin
      datar <= 16'b 1000001111010111;
      datai <= 16'b 0001111100011010;
      //552
    end
    10'b 1010111001 : begin
      datar <= 16'b 1000010001101111;
      datai <= 16'b 0010000101100001;
      //555
    end
    10'b 1010111010 : begin
      datar <= 16'b 1000010100010010;
      datai <= 16'b 0010001110100110;
      //558
    end
    10'b 1010111011 : begin
      datar <= 16'b 1000010110111111;
      datai <= 16'b 0010010111101000;
      //561
    end
    10'b 1010111100 : begin
      datar <= 16'b 1000011001110111;
      datai <= 16'b 0010100000100110;
      //564
    end
    10'b 1010111101 : begin
      datar <= 16'b 1000011100111001;
      datai <= 16'b 0010101001100001;
      //567
    end
    10'b 1010111110 : begin
      datar <= 16'b 1000100000000110;
      datai <= 16'b 0010110010011001;
      //570
    end
    10'b 1010111111 : begin
      datar <= 16'b 1000100011011110;
      datai <= 16'b 0010111011001100;
      //573
    end
    10'b 1011000000 : begin
      datar <= 16'b 1000100110111111;
      datai <= 16'b 0011000011111011;
      //576
    end
    10'b 1011000001 : begin
      datar <= 16'b 1000101010101011;
      datai <= 16'b 0011001100100110;
      //579
    end
    10'b 1011000010 : begin
      datar <= 16'b 1000101110100001;
      datai <= 16'b 0011010101001101;
      //582
    end
    10'b 1011000011 : begin
      datar <= 16'b 1000110010100010;
      datai <= 16'b 0011011101101111;
      //585
    end
    10'b 1011000100 : begin
      datar <= 16'b 1000110110101100;
      datai <= 16'b 0011100110001100;
      //588
    end
    10'b 1011000101 : begin
      datar <= 16'b 1000111011000000;
      datai <= 16'b 0011101110100101;
      //591
    end
    10'b 1011000110 : begin
      datar <= 16'b 1000111111011110;
      datai <= 16'b 0011110110111000;
      //594
    end
    10'b 1011000111 : begin
      datar <= 16'b 1001000100000101;
      datai <= 16'b 0011111111000101;
      //597
    end
    10'b 1011001000 : begin
      datar <= 16'b 1001001000110111;
      datai <= 16'b 0100000111001110;
      //600
    end
    10'b 1011001001 : begin
      datar <= 16'b 1001001101110010;
      datai <= 16'b 0100001111010000;
      //603
    end
    10'b 1011001010 : begin
      datar <= 16'b 1001010010110110;
      datai <= 16'b 0100010111001101;
      //606
    end
    10'b 1011001011 : begin
      datar <= 16'b 1001011000000011;
      datai <= 16'b 0100011111000011;
      //609
    end
    10'b 1011001100 : begin
      datar <= 16'b 1001011101011010;
      datai <= 16'b 0100100110110100;
      //612
    end
    10'b 1011001101 : begin
      datar <= 16'b 1001100010111010;
      datai <= 16'b 0100101110011101;
      //615
    end
    10'b 1011001110 : begin
      datar <= 16'b 1001101000100011;
      datai <= 16'b 0100110110000001;
      //618
    end
    10'b 1011001111 : begin
      datar <= 16'b 1001101110010100;
      datai <= 16'b 0100111101011101;
      //621
    end
    10'b 1011010000 : begin
      datar <= 16'b 1001110100001111;
      datai <= 16'b 0101000100110011;
      //624
    end
    10'b 1011010001 : begin
      datar <= 16'b 1001111010010010;
      datai <= 16'b 0101001100000010;
      //627
    end
    10'b 1011010010 : begin
      datar <= 16'b 1010000000011101;
      datai <= 16'b 0101010011001001;
      //630
    end
    10'b 1011010011 : begin
      datar <= 16'b 1010000110110001;
      datai <= 16'b 0101011010001010;
      //633
    end
    10'b 1011010100 : begin
      datar <= 16'b 1010001101001101;
      datai <= 16'b 0101100001000010;
      //636
    end
    10'b 1011010101 : begin
      datar <= 16'b 1010010011110001;
      datai <= 16'b 0101100111110011;
      //639
    end
    10'b 1011010110 : begin
      datar <= 16'b 1010011010011100;
      datai <= 16'b 0101101110011100;
      //642
    end
    10'b 1011010111 : begin
      datar <= 16'b 1010100001010000;
      datai <= 16'b 0101110100111110;
      //645
    end
    10'b 1011011000 : begin
      datar <= 16'b 1010101000001011;
      datai <= 16'b 0101111011010111;
      //648
    end
    10'b 1011011001 : begin
      datar <= 16'b 1010101111001110;
      datai <= 16'b 0110000001101000;
      //651
    end
    10'b 1011011010 : begin
      datar <= 16'b 1010110110011000;
      datai <= 16'b 0110000111110000;
      //654
    end
    10'b 1011011011 : begin
      datar <= 16'b 1010111101101001;
      datai <= 16'b 0110001101110000;
      //657
    end
    10'b 1011011100 : begin
      datar <= 16'b 1011000101000001;
      datai <= 16'b 0110010011101000;
      //660
    end
    10'b 1011011101 : begin
      datar <= 16'b 1011001100100000;
      datai <= 16'b 0110011001010110;
      //663
    end
    10'b 1011011110 : begin
      datar <= 16'b 1011010100000101;
      datai <= 16'b 0110011110111100;
      //666
    end
    10'b 1011011111 : begin
      datar <= 16'b 1011011011110001;
      datai <= 16'b 0110100100011001;
      //669
    end
    10'b 1011100000 : begin
      datar <= 16'b 1011100011100100;
      datai <= 16'b 0110101001101101;
      //672
    end
    10'b 1011100001 : begin
      datar <= 16'b 1011101011011100;
      datai <= 16'b 0110101110110111;
      //675
    end
    10'b 1011100010 : begin
      datar <= 16'b 1011110011011011;
      datai <= 16'b 0110110011111000;
      //678
    end
    10'b 1011100011 : begin
      datar <= 16'b 1011111011011111;
      datai <= 16'b 0110111000110000;
      //681
    end
    10'b 1011100100 : begin
      datar <= 16'b 1100000011101001;
      datai <= 16'b 0110111101011110;
      //684
    end
    10'b 1011100101 : begin
      datar <= 16'b 1100001011111001;
      datai <= 16'b 0111000010000011;
      //687
    end
    10'b 1011100110 : begin
      datar <= 16'b 1100010100001110;
      datai <= 16'b 0111000110011101;
      //690
    end
    10'b 1011100111 : begin
      datar <= 16'b 1100011100100111;
      datai <= 16'b 0111001010101110;
      //693
    end
    10'b 1011101000 : begin
      datar <= 16'b 1100100101000110;
      datai <= 16'b 0111001110110101;
      //696
    end
    10'b 1011101001 : begin
      datar <= 16'b 1100101101101010;
      datai <= 16'b 0111010010110010;
      //699
    end
    10'b 1011101010 : begin
      datar <= 16'b 1100110110010010;
      datai <= 16'b 0111010110100101;
      //702
    end
    10'b 1011101011 : begin
      datar <= 16'b 1100111110111111;
      datai <= 16'b 0111011010001101;
      //705
    end
    10'b 1011101100 : begin
      datar <= 16'b 1101000111101111;
      datai <= 16'b 0111011101101011;
      //708
    end
    10'b 1011101101 : begin
      datar <= 16'b 1101010000100100;
      datai <= 16'b 0111100000111111;
      //711
    end
    10'b 1011101110 : begin
      datar <= 16'b 1101011001011101;
      datai <= 16'b 0111100100001001;
      //714
    end
    10'b 1011101111 : begin
      datar <= 16'b 1101100010011001;
      datai <= 16'b 0111100111001000;
      //717
    end
    10'b 1011110000 : begin
      datar <= 16'b 1101101011011000;
      datai <= 16'b 0111101001111100;
      //720
    end
    10'b 1011110001 : begin
      datar <= 16'b 1101110100011011;
      datai <= 16'b 0111101100100110;
      //723
    end
    10'b 1011110010 : begin
      datar <= 16'b 1101111101100001;
      datai <= 16'b 0111101111000101;
      //726
    end
    10'b 1011110011 : begin
      datar <= 16'b 1110000110101001;
      datai <= 16'b 0111110001011001;
      //729
    end
    10'b 1011110100 : begin
      datar <= 16'b 1110001111110101;
      datai <= 16'b 0111110011100011;
      //732
    end
    10'b 1011110101 : begin
      datar <= 16'b 1110011001000010;
      datai <= 16'b 0111110101100010;
      //735
    end
    10'b 1011110110 : begin
      datar <= 16'b 1110100010010010;
      datai <= 16'b 0111110111010101;
      //738
    end
    10'b 1011110111 : begin
      datar <= 16'b 1110101011100100;
      datai <= 16'b 0111111000111110;
      //741
    end
    10'b 1011111000 : begin
      datar <= 16'b 1110110100111000;
      datai <= 16'b 0111111010011100;
      //744
    end
    10'b 1011111001 : begin
      datar <= 16'b 1110111110001110;
      datai <= 16'b 0111111011101111;
      //747
    end
    10'b 1011111010 : begin
      datar <= 16'b 1111000111100100;
      datai <= 16'b 0111111100110111;
      //750
    end
    10'b 1011111011 : begin
      datar <= 16'b 1111010000111100;
      datai <= 16'b 0111111101110100;
      //753
    end
    10'b 1011111100 : begin
      datar <= 16'b 1111011010010110;
      datai <= 16'b 0111111110100110;
      //756
    end
    10'b 1011111101 : begin
      datar <= 16'b 1111100011101111;
      datai <= 16'b 0111111111001101;
      //759
    end
    10'b 1011111110 : begin
      datar <= 16'b 1111101101001010;
      datai <= 16'b 0111111111101001;
      //762
    end
    10'b 1011111111 : begin
      datar <= 16'b 1111110110100101;
      datai <= 16'b 0111111111111001;
      //765
    end
    10'b 1100000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100000111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100001111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100010111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100011111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100100111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100101111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100110111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1100111111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101000111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101001111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101010111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101011111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101100111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101101111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101110111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1101111111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110000111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110001111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110010111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110011111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110100111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110101111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110110111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1110111111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111000111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111001111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111010111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111011111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111100111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111101111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111110111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    10'b 1111111111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    default : begin
      for (i=data_width - 1; i >= 0; i = i - 1) begin
        datar[i] <= 1'b 0;
        datai[i] <= 1'b 0;
      end
    end
    endcase
  end


endmodule
