// File ./rom2.vhd translated with vhd2vl v2.4 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 1995

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002, 2005, 2008-2010 Larry Doolittle - LBNL
//     http://doolittle.icarus.com/~larry/vhd2vl/
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

// Rom file for twiddle factors 
// ../../../rtl/vhdl/WISHBONE_FFT/rom2.vhd contains 256 points of 16 width 
//  for a 1024 point fft.
// no timescale needed

module rom2(
clk,
address,
datar,
datai
);

parameter [31:0] data_width=16;
parameter [31:0] address_width=8;
input clk;
input [7:0] address;
output [data_width - 1:0] datar;
output [data_width - 1:0] datai;

wire clk;
wire [7:0] address;
reg [data_width - 1:0] datar;
reg [data_width - 1:0] datai;
integer i;


  always @(posedge address or posedge clk) begin
    case(address)
    8'b 00000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 00000001 : begin
      datar <= 16'b 0111111111011000;
      datai <= 16'b 1111100110111000;
      //8
    end
    8'b 00000010 : begin
      datar <= 16'b 0111111101100001;
      datai <= 16'b 1111001101110100;
      //16
    end
    8'b 00000011 : begin
      datar <= 16'b 0111111010011100;
      datai <= 16'b 1110110100111000;
      //24
    end
    8'b 00000100 : begin
      datar <= 16'b 0111110110001001;
      datai <= 16'b 1110011100000111;
      //32
    end
    8'b 00000101 : begin
      datar <= 16'b 0111110000101001;
      datai <= 16'b 1110000011100110;
      //40
    end
    8'b 00000110 : begin
      datar <= 16'b 0111101001111100;
      datai <= 16'b 1101101011011000;
      //48
    end
    8'b 00000111 : begin
      datar <= 16'b 0111100010000100;
      datai <= 16'b 1101010011100001;
      //56
    end
    8'b 00001000 : begin
      datar <= 16'b 0111011001000001;
      datai <= 16'b 1100111100000101;
      //64
    end
    8'b 00001001 : begin
      datar <= 16'b 0111001110110101;
      datai <= 16'b 1100100101000110;
      //72
    end
    8'b 00001010 : begin
      datar <= 16'b 0111000011100010;
      datai <= 16'b 1100001110101010;
      //80
    end
    8'b 00001011 : begin
      datar <= 16'b 0110110111001001;
      datai <= 16'b 1011111000110010;
      //88
    end
    8'b 00001100 : begin
      datar <= 16'b 0110101001101101;
      datai <= 16'b 1011100011100100;
      //96
    end
    8'b 00001101 : begin
      datar <= 16'b 0110011011001111;
      datai <= 16'b 1011001111000001;
      //104
    end
    8'b 00001110 : begin
      datar <= 16'b 0110001011110001;
      datai <= 16'b 1010111011001101;
      //112
    end
    8'b 00001111 : begin
      datar <= 16'b 0101111011010111;
      datai <= 16'b 1010101000001011;
      //120
    end
    8'b 00010000 : begin
      datar <= 16'b 0101101010000010;
      datai <= 16'b 1010010101111110;
      //128
    end
    8'b 00010001 : begin
      datar <= 16'b 0101010111110101;
      datai <= 16'b 1010000100101001;
      //136
    end
    8'b 00010010 : begin
      datar <= 16'b 0101000100110011;
      datai <= 16'b 1001110100001111;
      //144
    end
    8'b 00010011 : begin
      datar <= 16'b 0100110000111111;
      datai <= 16'b 1001100100110001;
      //152
    end
    8'b 00010100 : begin
      datar <= 16'b 0100011100011100;
      datai <= 16'b 1001010110010011;
      //160
    end
    8'b 00010101 : begin
      datar <= 16'b 0100000111001110;
      datai <= 16'b 1001001000110111;
      //168
    end
    8'b 00010110 : begin
      datar <= 16'b 0011110001010110;
      datai <= 16'b 1000111100011110;
      //176
    end
    8'b 00010111 : begin
      datar <= 16'b 0011011010111010;
      datai <= 16'b 1000110001001011;
      //184
    end
    8'b 00011000 : begin
      datar <= 16'b 0011000011111011;
      datai <= 16'b 1000100110111111;
      //192
    end
    8'b 00011001 : begin
      datar <= 16'b 0010101100011111;
      datai <= 16'b 1000011101111100;
      //200
    end
    8'b 00011010 : begin
      datar <= 16'b 0010010100101000;
      datai <= 16'b 1000010110000100;
      //208
    end
    8'b 00011011 : begin
      datar <= 16'b 0001111100011010;
      datai <= 16'b 1000001111010111;
      //216
    end
    8'b 00011100 : begin
      datar <= 16'b 0001100011111001;
      datai <= 16'b 1000001001110111;
      //224
    end
    8'b 00011101 : begin
      datar <= 16'b 0001001011001000;
      datai <= 16'b 1000000101100100;
      //232
    end
    8'b 00011110 : begin
      datar <= 16'b 0000110010001100;
      datai <= 16'b 1000000010011111;
      //240
    end
    8'b 00011111 : begin
      datar <= 16'b 0000011001001000;
      datai <= 16'b 1000000000101000;
      //248
    end
    8'b 00100000 : begin
      datar <= 16'b 0000000000000000;
      datai <= 16'b 1000000000000001;
      //256
    end
    8'b 00100001 : begin
      datar <= 16'b 1111100110111000;
      datai <= 16'b 1000000000101000;
      //264
    end
    8'b 00100010 : begin
      datar <= 16'b 1111001101110100;
      datai <= 16'b 1000000010011111;
      //272
    end
    8'b 00100011 : begin
      datar <= 16'b 1110110100111000;
      datai <= 16'b 1000000101100100;
      //280
    end
    8'b 00100100 : begin
      datar <= 16'b 1110011100000111;
      datai <= 16'b 1000001001110111;
      //288
    end
    8'b 00100101 : begin
      datar <= 16'b 1110000011100110;
      datai <= 16'b 1000001111010111;
      //296
    end
    8'b 00100110 : begin
      datar <= 16'b 1101101011011000;
      datai <= 16'b 1000010110000100;
      //304
    end
    8'b 00100111 : begin
      datar <= 16'b 1101010011100001;
      datai <= 16'b 1000011101111100;
      //312
    end
    8'b 00101000 : begin
      datar <= 16'b 1100111100000101;
      datai <= 16'b 1000100110111111;
      //320
    end
    8'b 00101001 : begin
      datar <= 16'b 1100100101000110;
      datai <= 16'b 1000110001001011;
      //328
    end
    8'b 00101010 : begin
      datar <= 16'b 1100001110101010;
      datai <= 16'b 1000111100011110;
      //336
    end
    8'b 00101011 : begin
      datar <= 16'b 1011111000110010;
      datai <= 16'b 1001001000110111;
      //344
    end
    8'b 00101100 : begin
      datar <= 16'b 1011100011100100;
      datai <= 16'b 1001010110010011;
      //352
    end
    8'b 00101101 : begin
      datar <= 16'b 1011001111000001;
      datai <= 16'b 1001100100110001;
      //360
    end
    8'b 00101110 : begin
      datar <= 16'b 1010111011001101;
      datai <= 16'b 1001110100001111;
      //368
    end
    8'b 00101111 : begin
      datar <= 16'b 1010101000001011;
      datai <= 16'b 1010000100101001;
      //376
    end
    8'b 00110000 : begin
      datar <= 16'b 1010010101111110;
      datai <= 16'b 1010010101111110;
      //384
    end
    8'b 00110001 : begin
      datar <= 16'b 1010000100101001;
      datai <= 16'b 1010101000001011;
      //392
    end
    8'b 00110010 : begin
      datar <= 16'b 1001110100001111;
      datai <= 16'b 1010111011001101;
      //400
    end
    8'b 00110011 : begin
      datar <= 16'b 1001100100110001;
      datai <= 16'b 1011001111000001;
      //408
    end
    8'b 00110100 : begin
      datar <= 16'b 1001010110010011;
      datai <= 16'b 1011100011100100;
      //416
    end
    8'b 00110101 : begin
      datar <= 16'b 1001001000110111;
      datai <= 16'b 1011111000110010;
      //424
    end
    8'b 00110110 : begin
      datar <= 16'b 1000111100011110;
      datai <= 16'b 1100001110101010;
      //432
    end
    8'b 00110111 : begin
      datar <= 16'b 1000110001001011;
      datai <= 16'b 1100100101000110;
      //440
    end
    8'b 00111000 : begin
      datar <= 16'b 1000100110111111;
      datai <= 16'b 1100111100000101;
      //448
    end
    8'b 00111001 : begin
      datar <= 16'b 1000011101111100;
      datai <= 16'b 1101010011100001;
      //456
    end
    8'b 00111010 : begin
      datar <= 16'b 1000010110000100;
      datai <= 16'b 1101101011011000;
      //464
    end
    8'b 00111011 : begin
      datar <= 16'b 1000001111010111;
      datai <= 16'b 1110000011100110;
      //472
    end
    8'b 00111100 : begin
      datar <= 16'b 1000001001110111;
      datai <= 16'b 1110011100000111;
      //480
    end
    8'b 00111101 : begin
      datar <= 16'b 1000000101100100;
      datai <= 16'b 1110110100111000;
      //488
    end
    8'b 00111110 : begin
      datar <= 16'b 1000000010011111;
      datai <= 16'b 1111001101110100;
      //496
    end
    8'b 00111111 : begin
      datar <= 16'b 1000000000101000;
      datai <= 16'b 1111100110111000;
      //504
    end
    8'b 01000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 01000001 : begin
      datar <= 16'b 0111111111110101;
      datai <= 16'b 1111110011011100;
      //4
    end
    8'b 01000010 : begin
      datar <= 16'b 0111111111011000;
      datai <= 16'b 1111100110111000;
      //8
    end
    8'b 01000011 : begin
      datar <= 16'b 0111111110100110;
      datai <= 16'b 1111011010010110;
      //12
    end
    8'b 01000100 : begin
      datar <= 16'b 0111111101100001;
      datai <= 16'b 1111001101110100;
      //16
    end
    8'b 01000101 : begin
      datar <= 16'b 0111111100001001;
      datai <= 16'b 1111000001010101;
      //20
    end
    8'b 01000110 : begin
      datar <= 16'b 0111111010011100;
      datai <= 16'b 1110110100111000;
      //24
    end
    8'b 01000111 : begin
      datar <= 16'b 0111111000011101;
      datai <= 16'b 1110101000011110;
      //28
    end
    8'b 01001000 : begin
      datar <= 16'b 0111110110001001;
      datai <= 16'b 1110011100000111;
      //32
    end
    8'b 01001001 : begin
      datar <= 16'b 0111110011100011;
      datai <= 16'b 1110001111110101;
      //36
    end
    8'b 01001010 : begin
      datar <= 16'b 0111110000101001;
      datai <= 16'b 1110000011100110;
      //40
    end
    8'b 01001011 : begin
      datar <= 16'b 0111101101011100;
      datai <= 16'b 1101110111011101;
      //44
    end
    8'b 01001100 : begin
      datar <= 16'b 0111101001111100;
      datai <= 16'b 1101101011011000;
      //48
    end
    8'b 01001101 : begin
      datar <= 16'b 0111100110001001;
      datai <= 16'b 1101011111011010;
      //52
    end
    8'b 01001110 : begin
      datar <= 16'b 0111100010000100;
      datai <= 16'b 1101010011100001;
      //56
    end
    8'b 01001111 : begin
      datar <= 16'b 0111011101101011;
      datai <= 16'b 1101000111101111;
      //60
    end
    8'b 01010000 : begin
      datar <= 16'b 0111011001000001;
      datai <= 16'b 1100111100000101;
      //64
    end
    8'b 01010001 : begin
      datar <= 16'b 0111010100000100;
      datai <= 16'b 1100110000100001;
      //68
    end
    8'b 01010010 : begin
      datar <= 16'b 0111001110110101;
      datai <= 16'b 1100100101000110;
      //72
    end
    8'b 01010011 : begin
      datar <= 16'b 0111001001010100;
      datai <= 16'b 1100011001110100;
      //76
    end
    8'b 01010100 : begin
      datar <= 16'b 0111000011100010;
      datai <= 16'b 1100001110101010;
      //80
    end
    8'b 01010101 : begin
      datar <= 16'b 0110111101011110;
      datai <= 16'b 1100000011101001;
      //84
    end
    8'b 01010110 : begin
      datar <= 16'b 0110110111001001;
      datai <= 16'b 1011111000110010;
      //88
    end
    8'b 01010111 : begin
      datar <= 16'b 0110110000100011;
      datai <= 16'b 1011101110000110;
      //92
    end
    8'b 01011000 : begin
      datar <= 16'b 0110101001101101;
      datai <= 16'b 1011100011100100;
      //96
    end
    8'b 01011001 : begin
      datar <= 16'b 0110100010100110;
      datai <= 16'b 1011011001001100;
      //100
    end
    8'b 01011010 : begin
      datar <= 16'b 0110011011001111;
      datai <= 16'b 1011001111000001;
      //104
    end
    8'b 01011011 : begin
      datar <= 16'b 0110010011101000;
      datai <= 16'b 1011000101000001;
      //108
    end
    8'b 01011100 : begin
      datar <= 16'b 0110001011110001;
      datai <= 16'b 1010111011001101;
      //112
    end
    8'b 01011101 : begin
      datar <= 16'b 0110000011101011;
      datai <= 16'b 1010110001100101;
      //116
    end
    8'b 01011110 : begin
      datar <= 16'b 0101111011010111;
      datai <= 16'b 1010101000001011;
      //120
    end
    8'b 01011111 : begin
      datar <= 16'b 0101110010110011;
      datai <= 16'b 1010011110111110;
      //124
    end
    8'b 01100000 : begin
      datar <= 16'b 0101101010000010;
      datai <= 16'b 1010010101111110;
      //128
    end
    8'b 01100001 : begin
      datar <= 16'b 0101100001000010;
      datai <= 16'b 1010001101001101;
      //132
    end
    8'b 01100010 : begin
      datar <= 16'b 0101010111110101;
      datai <= 16'b 1010000100101001;
      //136
    end
    8'b 01100011 : begin
      datar <= 16'b 0101001110011011;
      datai <= 16'b 1001111100010101;
      //140
    end
    8'b 01100100 : begin
      datar <= 16'b 0101000100110011;
      datai <= 16'b 1001110100001111;
      //144
    end
    8'b 01100101 : begin
      datar <= 16'b 0100111010111111;
      datai <= 16'b 1001101100011000;
      //148
    end
    8'b 01100110 : begin
      datar <= 16'b 0100110000111111;
      datai <= 16'b 1001100100110001;
      //152
    end
    8'b 01100111 : begin
      datar <= 16'b 0100100110110100;
      datai <= 16'b 1001011101011010;
      //156
    end
    8'b 01101000 : begin
      datar <= 16'b 0100011100011100;
      datai <= 16'b 1001010110010011;
      //160
    end
    8'b 01101001 : begin
      datar <= 16'b 0100010001111010;
      datai <= 16'b 1001001111011101;
      //164
    end
    8'b 01101010 : begin
      datar <= 16'b 0100000111001110;
      datai <= 16'b 1001001000110111;
      //168
    end
    8'b 01101011 : begin
      datar <= 16'b 0011111100010111;
      datai <= 16'b 1001000010100010;
      //172
    end
    8'b 01101100 : begin
      datar <= 16'b 0011110001010110;
      datai <= 16'b 1000111100011110;
      //176
    end
    8'b 01101101 : begin
      datar <= 16'b 0011100110001100;
      datai <= 16'b 1000110110101100;
      //180
    end
    8'b 01101110 : begin
      datar <= 16'b 0011011010111010;
      datai <= 16'b 1000110001001011;
      //184
    end
    8'b 01101111 : begin
      datar <= 16'b 0011001111011111;
      datai <= 16'b 1000101011111100;
      //188
    end
    8'b 01110000 : begin
      datar <= 16'b 0011000011111011;
      datai <= 16'b 1000100110111111;
      //192
    end
    8'b 01110001 : begin
      datar <= 16'b 0010111000010001;
      datai <= 16'b 1000100010010101;
      //196
    end
    8'b 01110010 : begin
      datar <= 16'b 0010101100011111;
      datai <= 16'b 1000011101111100;
      //200
    end
    8'b 01110011 : begin
      datar <= 16'b 0010100000100110;
      datai <= 16'b 1000011001110111;
      //204
    end
    8'b 01110100 : begin
      datar <= 16'b 0010010100101000;
      datai <= 16'b 1000010110000100;
      //208
    end
    8'b 01110101 : begin
      datar <= 16'b 0010001000100011;
      datai <= 16'b 1000010010100100;
      //212
    end
    8'b 01110110 : begin
      datar <= 16'b 0001111100011010;
      datai <= 16'b 1000001111010111;
      //216
    end
    8'b 01110111 : begin
      datar <= 16'b 0001110000001011;
      datai <= 16'b 1000001100011101;
      //220
    end
    8'b 01111000 : begin
      datar <= 16'b 0001100011111001;
      datai <= 16'b 1000001001110111;
      //224
    end
    8'b 01111001 : begin
      datar <= 16'b 0001010111100010;
      datai <= 16'b 1000000111100011;
      //228
    end
    8'b 01111010 : begin
      datar <= 16'b 0001001011001000;
      datai <= 16'b 1000000101100100;
      //232
    end
    8'b 01111011 : begin
      datar <= 16'b 0000111110101011;
      datai <= 16'b 1000000011110111;
      //236
    end
    8'b 01111100 : begin
      datar <= 16'b 0000110010001100;
      datai <= 16'b 1000000010011111;
      //240
    end
    8'b 01111101 : begin
      datar <= 16'b 0000100101101010;
      datai <= 16'b 1000000001011010;
      //244
    end
    8'b 01111110 : begin
      datar <= 16'b 0000011001001000;
      datai <= 16'b 1000000000101000;
      //248
    end
    8'b 01111111 : begin
      datar <= 16'b 0000001100100100;
      datai <= 16'b 1000000000001011;
      //252
    end
    8'b 10000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 10000001 : begin
      datar <= 16'b 0111111110100110;
      datai <= 16'b 1111011010010110;
      //12
    end
    8'b 10000010 : begin
      datar <= 16'b 0111111010011100;
      datai <= 16'b 1110110100111000;
      //24
    end
    8'b 10000011 : begin
      datar <= 16'b 0111110011100011;
      datai <= 16'b 1110001111110101;
      //36
    end
    8'b 10000100 : begin
      datar <= 16'b 0111101001111100;
      datai <= 16'b 1101101011011000;
      //48
    end
    8'b 10000101 : begin
      datar <= 16'b 0111011101101011;
      datai <= 16'b 1101000111101111;
      //60
    end
    8'b 10000110 : begin
      datar <= 16'b 0111001110110101;
      datai <= 16'b 1100100101000110;
      //72
    end
    8'b 10000111 : begin
      datar <= 16'b 0110111101011110;
      datai <= 16'b 1100000011101001;
      //84
    end
    8'b 10001000 : begin
      datar <= 16'b 0110101001101101;
      datai <= 16'b 1011100011100100;
      //96
    end
    8'b 10001001 : begin
      datar <= 16'b 0110010011101000;
      datai <= 16'b 1011000101000001;
      //108
    end
    8'b 10001010 : begin
      datar <= 16'b 0101111011010111;
      datai <= 16'b 1010101000001011;
      //120
    end
    8'b 10001011 : begin
      datar <= 16'b 0101100001000010;
      datai <= 16'b 1010001101001101;
      //132
    end
    8'b 10001100 : begin
      datar <= 16'b 0101000100110011;
      datai <= 16'b 1001110100001111;
      //144
    end
    8'b 10001101 : begin
      datar <= 16'b 0100100110110100;
      datai <= 16'b 1001011101011010;
      //156
    end
    8'b 10001110 : begin
      datar <= 16'b 0100000111001110;
      datai <= 16'b 1001001000110111;
      //168
    end
    8'b 10001111 : begin
      datar <= 16'b 0011100110001100;
      datai <= 16'b 1000110110101100;
      //180
    end
    8'b 10010000 : begin
      datar <= 16'b 0011000011111011;
      datai <= 16'b 1000100110111111;
      //192
    end
    8'b 10010001 : begin
      datar <= 16'b 0010100000100110;
      datai <= 16'b 1000011001110111;
      //204
    end
    8'b 10010010 : begin
      datar <= 16'b 0001111100011010;
      datai <= 16'b 1000001111010111;
      //216
    end
    8'b 10010011 : begin
      datar <= 16'b 0001010111100010;
      datai <= 16'b 1000000111100011;
      //228
    end
    8'b 10010100 : begin
      datar <= 16'b 0000110010001100;
      datai <= 16'b 1000000010011111;
      //240
    end
    8'b 10010101 : begin
      datar <= 16'b 0000001100100100;
      datai <= 16'b 1000000000001011;
      //252
    end
    8'b 10010110 : begin
      datar <= 16'b 1111100110111000;
      datai <= 16'b 1000000000101000;
      //264
    end
    8'b 10010111 : begin
      datar <= 16'b 1111000001010101;
      datai <= 16'b 1000000011110111;
      //276
    end
    8'b 10011000 : begin
      datar <= 16'b 1110011100000111;
      datai <= 16'b 1000001001110111;
      //288
    end
    8'b 10011001 : begin
      datar <= 16'b 1101110111011101;
      datai <= 16'b 1000010010100100;
      //300
    end
    8'b 10011010 : begin
      datar <= 16'b 1101010011100001;
      datai <= 16'b 1000011101111100;
      //312
    end
    8'b 10011011 : begin
      datar <= 16'b 1100110000100001;
      datai <= 16'b 1000101011111100;
      //324
    end
    8'b 10011100 : begin
      datar <= 16'b 1100001110101010;
      datai <= 16'b 1000111100011110;
      //336
    end
    8'b 10011101 : begin
      datar <= 16'b 1011101110000110;
      datai <= 16'b 1001001111011101;
      //348
    end
    8'b 10011110 : begin
      datar <= 16'b 1011001111000001;
      datai <= 16'b 1001100100110001;
      //360
    end
    8'b 10011111 : begin
      datar <= 16'b 1010110001100101;
      datai <= 16'b 1001111100010101;
      //372
    end
    8'b 10100000 : begin
      datar <= 16'b 1010010101111110;
      datai <= 16'b 1010010101111110;
      //384
    end
    8'b 10100001 : begin
      datar <= 16'b 1001111100010101;
      datai <= 16'b 1010110001100101;
      //396
    end
    8'b 10100010 : begin
      datar <= 16'b 1001100100110001;
      datai <= 16'b 1011001111000001;
      //408
    end
    8'b 10100011 : begin
      datar <= 16'b 1001001111011101;
      datai <= 16'b 1011101110000110;
      //420
    end
    8'b 10100100 : begin
      datar <= 16'b 1000111100011110;
      datai <= 16'b 1100001110101010;
      //432
    end
    8'b 10100101 : begin
      datar <= 16'b 1000101011111100;
      datai <= 16'b 1100110000100001;
      //444
    end
    8'b 10100110 : begin
      datar <= 16'b 1000011101111100;
      datai <= 16'b 1101010011100001;
      //456
    end
    8'b 10100111 : begin
      datar <= 16'b 1000010010100100;
      datai <= 16'b 1101110111011101;
      //468
    end
    8'b 10101000 : begin
      datar <= 16'b 1000001001110111;
      datai <= 16'b 1110011100000111;
      //480
    end
    8'b 10101001 : begin
      datar <= 16'b 1000000011110111;
      datai <= 16'b 1111000001010101;
      //492
    end
    8'b 10101010 : begin
      datar <= 16'b 1000000000101000;
      datai <= 16'b 1111100110111000;
      //504
    end
    8'b 10101011 : begin
      datar <= 16'b 1000000000001011;
      datai <= 16'b 0000001100100100;
      //516
    end
    8'b 10101100 : begin
      datar <= 16'b 1000000010011111;
      datai <= 16'b 0000110010001100;
      //528
    end
    8'b 10101101 : begin
      datar <= 16'b 1000000111100011;
      datai <= 16'b 0001010111100010;
      //540
    end
    8'b 10101110 : begin
      datar <= 16'b 1000001111010111;
      datai <= 16'b 0001111100011010;
      //552
    end
    8'b 10101111 : begin
      datar <= 16'b 1000011001110111;
      datai <= 16'b 0010100000100110;
      //564
    end
    8'b 10110000 : begin
      datar <= 16'b 1000100110111111;
      datai <= 16'b 0011000011111011;
      //576
    end
    8'b 10110001 : begin
      datar <= 16'b 1000110110101100;
      datai <= 16'b 0011100110001100;
      //588
    end
    8'b 10110010 : begin
      datar <= 16'b 1001001000110111;
      datai <= 16'b 0100000111001110;
      //600
    end
    8'b 10110011 : begin
      datar <= 16'b 1001011101011010;
      datai <= 16'b 0100100110110100;
      //612
    end
    8'b 10110100 : begin
      datar <= 16'b 1001110100001111;
      datai <= 16'b 0101000100110011;
      //624
    end
    8'b 10110101 : begin
      datar <= 16'b 1010001101001101;
      datai <= 16'b 0101100001000010;
      //636
    end
    8'b 10110110 : begin
      datar <= 16'b 1010101000001011;
      datai <= 16'b 0101111011010111;
      //648
    end
    8'b 10110111 : begin
      datar <= 16'b 1011000101000001;
      datai <= 16'b 0110010011101000;
      //660
    end
    8'b 10111000 : begin
      datar <= 16'b 1011100011100100;
      datai <= 16'b 0110101001101101;
      //672
    end
    8'b 10111001 : begin
      datar <= 16'b 1100000011101001;
      datai <= 16'b 0110111101011110;
      //684
    end
    8'b 10111010 : begin
      datar <= 16'b 1100100101000110;
      datai <= 16'b 0111001110110101;
      //696
    end
    8'b 10111011 : begin
      datar <= 16'b 1101000111101111;
      datai <= 16'b 0111011101101011;
      //708
    end
    8'b 10111100 : begin
      datar <= 16'b 1101101011011000;
      datai <= 16'b 0111101001111100;
      //720
    end
    8'b 10111101 : begin
      datar <= 16'b 1110001111110101;
      datai <= 16'b 0111110011100011;
      //732
    end
    8'b 10111110 : begin
      datar <= 16'b 1110110100111000;
      datai <= 16'b 0111111010011100;
      //744
    end
    8'b 10111111 : begin
      datar <= 16'b 1111011010010110;
      datai <= 16'b 0111111110100110;
      //756
    end
    8'b 11000000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11000111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11001111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11010111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11011111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11100111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11101111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11110111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111000 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111001 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111010 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111011 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111100 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111101 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111110 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    8'b 11111111 : begin
      datar <= 16'b 0111111111111111;
      datai <= 16'b 0000000000000000;
      //0
    end
    default : begin
      for (i=data_width - 1; i >= 0; i = i - 1) begin
        datar[i] <= 1'b 0;
        datai[i] <= 1'b 0;
      end
    end
    endcase
  end


endmodule
